module tt_um_cattuto_sr_latch (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input VPWR;
 input VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \shift_reg[0].genblk1.latch.clk ;
 wire \shift_reg[0].genblk1.latch.q ;
 wire \shift_reg[100].genblk1.genblk1.latch.clk ;
 wire \shift_reg[100].genblk1.genblk1.latch.clkout ;
 wire \shift_reg[100].genblk1.genblk1.latch.d ;
 wire \shift_reg[100].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[100].genblk1.genblk1.latch.q ;
 wire \shift_reg[101].genblk1.genblk1.latch.clk ;
 wire \shift_reg[101].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[101].genblk1.genblk1.latch.q ;
 wire \shift_reg[102].genblk1.genblk1.latch.clk ;
 wire \shift_reg[102].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[102].genblk1.genblk1.latch.q ;
 wire \shift_reg[103].genblk1.genblk1.latch.clk ;
 wire \shift_reg[103].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[103].genblk1.genblk1.latch.q ;
 wire \shift_reg[104].genblk1.genblk1.latch.clk ;
 wire \shift_reg[104].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[104].genblk1.genblk1.latch.q ;
 wire \shift_reg[105].genblk1.genblk1.latch.clk ;
 wire \shift_reg[105].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[105].genblk1.genblk1.latch.q ;
 wire \shift_reg[106].genblk1.genblk1.latch.clk ;
 wire \shift_reg[106].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[106].genblk1.genblk1.latch.q ;
 wire \shift_reg[107].genblk1.genblk1.latch.clk ;
 wire \shift_reg[107].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[107].genblk1.genblk1.latch.q ;
 wire \shift_reg[108].genblk1.genblk1.latch.clk ;
 wire \shift_reg[108].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[108].genblk1.genblk1.latch.q ;
 wire \shift_reg[109].genblk1.genblk1.latch.clk ;
 wire \shift_reg[109].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[109].genblk1.genblk1.latch.q ;
 wire \shift_reg[10].genblk1.genblk1.latch.clk ;
 wire \shift_reg[10].genblk1.genblk1.latch.clkout ;
 wire \shift_reg[10].genblk1.genblk1.latch.d ;
 wire \shift_reg[10].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[10].genblk1.genblk1.latch.q ;
 wire \shift_reg[110].genblk1.genblk1.latch.clk ;
 wire \shift_reg[110].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[110].genblk1.genblk1.latch.q ;
 wire \shift_reg[111].genblk1.genblk1.latch.clk ;
 wire \shift_reg[111].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[111].genblk1.genblk1.latch.q ;
 wire \shift_reg[112].genblk1.genblk1.latch.clk ;
 wire \shift_reg[112].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[112].genblk1.genblk1.latch.q ;
 wire \shift_reg[113].genblk1.genblk1.latch.clk ;
 wire \shift_reg[113].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[113].genblk1.genblk1.latch.q ;
 wire \shift_reg[114].genblk1.genblk1.latch.clk ;
 wire \shift_reg[114].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[114].genblk1.genblk1.latch.q ;
 wire \shift_reg[115].genblk1.genblk1.latch.clk ;
 wire \shift_reg[115].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[115].genblk1.genblk1.latch.q ;
 wire \shift_reg[116].genblk1.genblk1.latch.clk ;
 wire \shift_reg[116].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[116].genblk1.genblk1.latch.q ;
 wire \shift_reg[117].genblk1.genblk1.latch.clk ;
 wire \shift_reg[117].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[117].genblk1.genblk1.latch.q ;
 wire \shift_reg[118].genblk1.genblk1.latch.clk ;
 wire \shift_reg[118].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[118].genblk1.genblk1.latch.q ;
 wire \shift_reg[119].genblk1.genblk1.latch.clk ;
 wire \shift_reg[119].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[119].genblk1.genblk1.latch.q ;
 wire \shift_reg[11].genblk1.genblk1.latch.clk ;
 wire \shift_reg[11].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[11].genblk1.genblk1.latch.q ;
 wire \shift_reg[120].genblk1.genblk1.latch.clk ;
 wire \shift_reg[120].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[120].genblk1.genblk1.latch.q ;
 wire \shift_reg[121].genblk1.genblk1.latch.clk ;
 wire \shift_reg[121].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[121].genblk1.genblk1.latch.q ;
 wire \shift_reg[122].genblk1.genblk1.latch.clk ;
 wire \shift_reg[122].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[122].genblk1.genblk1.latch.q ;
 wire \shift_reg[123].genblk1.genblk1.latch.clk ;
 wire \shift_reg[123].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[123].genblk1.genblk1.latch.q ;
 wire \shift_reg[124].genblk1.genblk1.latch.clk ;
 wire \shift_reg[124].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[124].genblk1.genblk1.latch.q ;
 wire \shift_reg[125].genblk1.genblk1.latch.clk ;
 wire \shift_reg[125].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[125].genblk1.genblk1.latch.q ;
 wire \shift_reg[126].genblk1.genblk1.latch.clk ;
 wire \shift_reg[126].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[126].genblk1.genblk1.latch.q ;
 wire \shift_reg[127].genblk1.genblk1.latch.clk ;
 wire \shift_reg[127].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[127].genblk1.genblk1.latch.q ;
 wire \shift_reg[128].genblk1.genblk1.latch.clk ;
 wire \shift_reg[128].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[128].genblk1.genblk1.latch.q ;
 wire \shift_reg[129].genblk1.genblk1.latch.clk ;
 wire \shift_reg[129].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[129].genblk1.genblk1.latch.q ;
 wire \shift_reg[12].genblk1.genblk1.latch.clk ;
 wire \shift_reg[12].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[12].genblk1.genblk1.latch.q ;
 wire \shift_reg[130].genblk1.genblk1.latch.clk ;
 wire \shift_reg[130].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[130].genblk1.genblk1.latch.q ;
 wire \shift_reg[131].genblk1.genblk1.latch.clk ;
 wire \shift_reg[131].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[131].genblk1.genblk1.latch.q ;
 wire \shift_reg[132].genblk1.genblk1.latch.clk ;
 wire \shift_reg[132].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[132].genblk1.genblk1.latch.q ;
 wire \shift_reg[133].genblk1.genblk1.latch.clk ;
 wire \shift_reg[133].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[133].genblk1.genblk1.latch.q ;
 wire \shift_reg[134].genblk1.genblk1.latch.clk ;
 wire \shift_reg[134].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[134].genblk1.genblk1.latch.q ;
 wire \shift_reg[135].genblk1.genblk1.latch.clk ;
 wire \shift_reg[135].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[135].genblk1.genblk1.latch.q ;
 wire \shift_reg[136].genblk1.genblk1.latch.clk ;
 wire \shift_reg[136].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[136].genblk1.genblk1.latch.q ;
 wire \shift_reg[137].genblk1.genblk1.latch.clk ;
 wire \shift_reg[137].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[137].genblk1.genblk1.latch.q ;
 wire \shift_reg[138].genblk1.genblk1.latch.clk ;
 wire \shift_reg[138].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[138].genblk1.genblk1.latch.q ;
 wire \shift_reg[139].genblk1.genblk1.latch.clk ;
 wire \shift_reg[139].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[139].genblk1.genblk1.latch.q ;
 wire \shift_reg[13].genblk1.genblk1.latch.clk ;
 wire \shift_reg[13].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[13].genblk1.genblk1.latch.q ;
 wire \shift_reg[140].genblk1.genblk1.latch.clk ;
 wire \shift_reg[140].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[140].genblk1.genblk1.latch.q ;
 wire \shift_reg[141].genblk1.genblk1.latch.clk ;
 wire \shift_reg[141].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[141].genblk1.genblk1.latch.q ;
 wire \shift_reg[142].genblk1.genblk1.latch.clk ;
 wire \shift_reg[142].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[142].genblk1.genblk1.latch.q ;
 wire \shift_reg[143].genblk1.genblk1.latch.clk ;
 wire \shift_reg[143].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[143].genblk1.genblk1.latch.q ;
 wire \shift_reg[144].genblk1.genblk1.latch.clk ;
 wire \shift_reg[144].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[144].genblk1.genblk1.latch.q ;
 wire \shift_reg[145].genblk1.genblk1.latch.clk ;
 wire \shift_reg[145].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[145].genblk1.genblk1.latch.q ;
 wire \shift_reg[146].genblk1.genblk1.latch.clk ;
 wire \shift_reg[146].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[146].genblk1.genblk1.latch.q ;
 wire \shift_reg[147].genblk1.genblk1.latch.clk ;
 wire \shift_reg[147].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[147].genblk1.genblk1.latch.q ;
 wire \shift_reg[148].genblk1.genblk1.latch.clk ;
 wire \shift_reg[148].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[148].genblk1.genblk1.latch.q ;
 wire \shift_reg[149].genblk1.genblk1.latch.clk ;
 wire \shift_reg[149].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[149].genblk1.genblk1.latch.q ;
 wire \shift_reg[14].genblk1.genblk1.latch.clk ;
 wire \shift_reg[14].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[14].genblk1.genblk1.latch.q ;
 wire \shift_reg[150].genblk1.genblk1.latch.clk ;
 wire \shift_reg[150].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[150].genblk1.genblk1.latch.q ;
 wire \shift_reg[151].genblk1.genblk1.latch.clk ;
 wire \shift_reg[151].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[151].genblk1.genblk1.latch.q ;
 wire \shift_reg[152].genblk1.genblk1.latch.clk ;
 wire \shift_reg[152].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[152].genblk1.genblk1.latch.q ;
 wire \shift_reg[153].genblk1.genblk1.latch.clk ;
 wire \shift_reg[153].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[153].genblk1.genblk1.latch.q ;
 wire \shift_reg[154].genblk1.genblk1.latch.clk ;
 wire \shift_reg[154].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[154].genblk1.genblk1.latch.q ;
 wire \shift_reg[155].genblk1.genblk1.latch.clk ;
 wire \shift_reg[155].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[155].genblk1.genblk1.latch.q ;
 wire \shift_reg[156].genblk1.genblk1.latch.clk ;
 wire \shift_reg[156].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[156].genblk1.genblk1.latch.q ;
 wire \shift_reg[157].genblk1.genblk1.latch.clk ;
 wire \shift_reg[157].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[157].genblk1.genblk1.latch.q ;
 wire \shift_reg[158].genblk1.genblk1.latch.clk ;
 wire \shift_reg[158].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[158].genblk1.genblk1.latch.q ;
 wire \shift_reg[159].genblk1.genblk1.latch.clk ;
 wire \shift_reg[159].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[159].genblk1.genblk1.latch.q ;
 wire \shift_reg[15].genblk1.genblk1.latch.clk ;
 wire \shift_reg[15].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[15].genblk1.genblk1.latch.q ;
 wire \shift_reg[160].genblk1.genblk1.latch.clk ;
 wire \shift_reg[160].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[160].genblk1.genblk1.latch.q ;
 wire \shift_reg[161].genblk1.genblk1.latch.clk ;
 wire \shift_reg[161].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[161].genblk1.genblk1.latch.q ;
 wire \shift_reg[162].genblk1.genblk1.latch.clk ;
 wire \shift_reg[162].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[162].genblk1.genblk1.latch.q ;
 wire \shift_reg[163].genblk1.genblk1.latch.clk ;
 wire \shift_reg[163].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[163].genblk1.genblk1.latch.q ;
 wire \shift_reg[164].genblk1.genblk1.latch.clk ;
 wire \shift_reg[164].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[164].genblk1.genblk1.latch.q ;
 wire \shift_reg[165].genblk1.genblk1.latch.clk ;
 wire \shift_reg[165].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[165].genblk1.genblk1.latch.q ;
 wire \shift_reg[166].genblk1.genblk1.latch.clk ;
 wire \shift_reg[166].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[166].genblk1.genblk1.latch.q ;
 wire \shift_reg[167].genblk1.genblk1.latch.clk ;
 wire \shift_reg[167].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[167].genblk1.genblk1.latch.q ;
 wire \shift_reg[168].genblk1.genblk1.latch.clk ;
 wire \shift_reg[168].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[168].genblk1.genblk1.latch.q ;
 wire \shift_reg[169].genblk1.genblk1.latch.clk ;
 wire \shift_reg[169].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[169].genblk1.genblk1.latch.q ;
 wire \shift_reg[16].genblk1.genblk1.latch.clk ;
 wire \shift_reg[16].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[16].genblk1.genblk1.latch.q ;
 wire \shift_reg[170].genblk1.genblk1.latch.clk ;
 wire \shift_reg[170].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[170].genblk1.genblk1.latch.q ;
 wire \shift_reg[171].genblk1.genblk1.latch.clk ;
 wire \shift_reg[171].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[171].genblk1.genblk1.latch.q ;
 wire \shift_reg[172].genblk1.genblk1.latch.clk ;
 wire \shift_reg[172].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[172].genblk1.genblk1.latch.q ;
 wire \shift_reg[173].genblk1.genblk1.latch.clk ;
 wire \shift_reg[173].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[173].genblk1.genblk1.latch.q ;
 wire \shift_reg[174].genblk1.genblk1.latch.clk ;
 wire \shift_reg[174].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[174].genblk1.genblk1.latch.q ;
 wire \shift_reg[175].genblk1.genblk1.latch.clk ;
 wire \shift_reg[175].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[175].genblk1.genblk1.latch.q ;
 wire \shift_reg[176].genblk1.genblk1.latch.clk ;
 wire \shift_reg[176].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[176].genblk1.genblk1.latch.q ;
 wire \shift_reg[177].genblk1.genblk1.latch.clk ;
 wire \shift_reg[177].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[177].genblk1.genblk1.latch.q ;
 wire \shift_reg[178].genblk1.genblk1.latch.clk ;
 wire \shift_reg[178].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[178].genblk1.genblk1.latch.q ;
 wire \shift_reg[179].genblk1.genblk1.latch.clk ;
 wire \shift_reg[179].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[179].genblk1.genblk1.latch.q ;
 wire \shift_reg[17].genblk1.genblk1.latch.clk ;
 wire \shift_reg[17].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[17].genblk1.genblk1.latch.q ;
 wire \shift_reg[180].genblk1.genblk1.latch.clk ;
 wire \shift_reg[180].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[180].genblk1.genblk1.latch.q ;
 wire \shift_reg[181].genblk1.genblk1.latch.clk ;
 wire \shift_reg[181].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[181].genblk1.genblk1.latch.q ;
 wire \shift_reg[182].genblk1.genblk1.latch.clk ;
 wire \shift_reg[182].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[182].genblk1.genblk1.latch.q ;
 wire \shift_reg[183].genblk1.genblk1.latch.clk ;
 wire \shift_reg[183].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[183].genblk1.genblk1.latch.q ;
 wire \shift_reg[184].genblk1.genblk1.latch.clk ;
 wire \shift_reg[184].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[184].genblk1.genblk1.latch.q ;
 wire \shift_reg[185].genblk1.genblk1.latch.clk ;
 wire \shift_reg[185].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[185].genblk1.genblk1.latch.q ;
 wire \shift_reg[186].genblk1.genblk1.latch.clk ;
 wire \shift_reg[186].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[186].genblk1.genblk1.latch.q ;
 wire \shift_reg[187].genblk1.genblk1.latch.clk ;
 wire \shift_reg[187].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[187].genblk1.genblk1.latch.q ;
 wire \shift_reg[188].genblk1.genblk1.latch.clk ;
 wire \shift_reg[188].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[188].genblk1.genblk1.latch.q ;
 wire \shift_reg[189].genblk1.genblk1.latch.clk ;
 wire \shift_reg[189].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[189].genblk1.genblk1.latch.q ;
 wire \shift_reg[18].genblk1.genblk1.latch.clk ;
 wire \shift_reg[18].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[18].genblk1.genblk1.latch.q ;
 wire \shift_reg[190].genblk1.genblk1.latch.clk ;
 wire \shift_reg[190].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[190].genblk1.genblk1.latch.q ;
 wire \shift_reg[191].genblk1.genblk1.latch.clk ;
 wire \shift_reg[191].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[191].genblk1.genblk1.latch.q ;
 wire \shift_reg[192].genblk1.genblk1.latch.clk ;
 wire \shift_reg[192].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[192].genblk1.genblk1.latch.q ;
 wire \shift_reg[193].genblk1.genblk1.latch.clk ;
 wire \shift_reg[193].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[193].genblk1.genblk1.latch.q ;
 wire \shift_reg[194].genblk1.genblk1.latch.clk ;
 wire \shift_reg[194].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[194].genblk1.genblk1.latch.q ;
 wire \shift_reg[195].genblk1.genblk1.latch.clk ;
 wire \shift_reg[195].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[195].genblk1.genblk1.latch.q ;
 wire \shift_reg[196].genblk1.genblk1.latch.clk ;
 wire \shift_reg[196].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[196].genblk1.genblk1.latch.q ;
 wire \shift_reg[197].genblk1.genblk1.latch.clk ;
 wire \shift_reg[197].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[197].genblk1.genblk1.latch.q ;
 wire \shift_reg[198].genblk1.genblk1.latch.clk ;
 wire \shift_reg[198].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[198].genblk1.genblk1.latch.q ;
 wire \shift_reg[199].genblk1.genblk1.latch.clk ;
 wire \shift_reg[199].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[199].genblk1.genblk1.latch.q ;
 wire \shift_reg[19].genblk1.genblk1.latch.clk ;
 wire \shift_reg[19].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[19].genblk1.genblk1.latch.q ;
 wire \shift_reg[1].genblk1.genblk1.latch.clk ;
 wire \shift_reg[1].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[1].genblk1.genblk1.latch.q ;
 wire \shift_reg[200].genblk1.genblk1.latch.clk ;
 wire \shift_reg[200].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[200].genblk1.genblk1.latch.q ;
 wire \shift_reg[201].genblk1.genblk1.latch.clk ;
 wire \shift_reg[201].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[201].genblk1.genblk1.latch.q ;
 wire \shift_reg[202].genblk1.genblk1.latch.clk ;
 wire \shift_reg[202].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[202].genblk1.genblk1.latch.q ;
 wire \shift_reg[203].genblk1.genblk1.latch.clk ;
 wire \shift_reg[203].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[203].genblk1.genblk1.latch.q ;
 wire \shift_reg[204].genblk1.genblk1.latch.clk ;
 wire \shift_reg[204].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[204].genblk1.genblk1.latch.q ;
 wire \shift_reg[205].genblk1.genblk1.latch.clk ;
 wire \shift_reg[205].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[205].genblk1.genblk1.latch.q ;
 wire \shift_reg[206].genblk1.genblk1.latch.clk ;
 wire \shift_reg[206].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[206].genblk1.genblk1.latch.q ;
 wire \shift_reg[207].genblk1.genblk1.latch.clk ;
 wire \shift_reg[207].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[207].genblk1.genblk1.latch.q ;
 wire \shift_reg[208].genblk1.genblk1.latch.clk ;
 wire \shift_reg[208].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[208].genblk1.genblk1.latch.q ;
 wire \shift_reg[209].genblk1.genblk1.latch.clk ;
 wire \shift_reg[209].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[209].genblk1.genblk1.latch.q ;
 wire \shift_reg[20].genblk1.genblk1.latch.clk ;
 wire \shift_reg[20].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[20].genblk1.genblk1.latch.q ;
 wire \shift_reg[210].genblk1.genblk1.latch.clk ;
 wire \shift_reg[210].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[210].genblk1.genblk1.latch.q ;
 wire \shift_reg[211].genblk1.genblk1.latch.clk ;
 wire \shift_reg[211].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[211].genblk1.genblk1.latch.q ;
 wire \shift_reg[212].genblk1.genblk1.latch.clk ;
 wire \shift_reg[212].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[212].genblk1.genblk1.latch.q ;
 wire \shift_reg[213].genblk1.genblk1.latch.clk ;
 wire \shift_reg[213].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[213].genblk1.genblk1.latch.q ;
 wire \shift_reg[214].genblk1.genblk1.latch.clk ;
 wire \shift_reg[214].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[214].genblk1.genblk1.latch.q ;
 wire \shift_reg[215].genblk1.genblk1.latch.clk ;
 wire \shift_reg[215].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[215].genblk1.genblk1.latch.q ;
 wire \shift_reg[216].genblk1.genblk1.latch.clk ;
 wire \shift_reg[216].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[216].genblk1.genblk1.latch.q ;
 wire \shift_reg[217].genblk1.genblk1.latch.clk ;
 wire \shift_reg[217].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[217].genblk1.genblk1.latch.q ;
 wire \shift_reg[218].genblk1.genblk1.latch.clk ;
 wire \shift_reg[218].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[218].genblk1.genblk1.latch.q ;
 wire \shift_reg[219].genblk1.genblk1.latch.clk ;
 wire \shift_reg[219].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[219].genblk1.genblk1.latch.q ;
 wire \shift_reg[21].genblk1.genblk1.latch.clk ;
 wire \shift_reg[21].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[21].genblk1.genblk1.latch.q ;
 wire \shift_reg[220].genblk1.genblk1.latch.clk ;
 wire \shift_reg[220].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[220].genblk1.genblk1.latch.q ;
 wire \shift_reg[221].genblk1.genblk1.latch.clk ;
 wire \shift_reg[221].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[221].genblk1.genblk1.latch.q ;
 wire \shift_reg[222].genblk1.genblk1.latch.clk ;
 wire \shift_reg[222].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[222].genblk1.genblk1.latch.q ;
 wire \shift_reg[223].genblk1.genblk1.latch.clk ;
 wire \shift_reg[223].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[223].genblk1.genblk1.latch.q ;
 wire \shift_reg[224].genblk1.genblk1.latch.clk ;
 wire \shift_reg[224].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[224].genblk1.genblk1.latch.q ;
 wire \shift_reg[225].genblk1.genblk1.latch.clk ;
 wire \shift_reg[225].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[225].genblk1.genblk1.latch.q ;
 wire \shift_reg[226].genblk1.genblk1.latch.clk ;
 wire \shift_reg[226].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[226].genblk1.genblk1.latch.q ;
 wire \shift_reg[227].genblk1.genblk1.latch.clk ;
 wire \shift_reg[227].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[227].genblk1.genblk1.latch.q ;
 wire \shift_reg[228].genblk1.genblk1.latch.clk ;
 wire \shift_reg[228].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[228].genblk1.genblk1.latch.q ;
 wire \shift_reg[229].genblk1.genblk1.latch.clk ;
 wire \shift_reg[229].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[229].genblk1.genblk1.latch.q ;
 wire \shift_reg[22].genblk1.genblk1.latch.clk ;
 wire \shift_reg[22].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[22].genblk1.genblk1.latch.q ;
 wire \shift_reg[230].genblk1.genblk1.latch.clk ;
 wire \shift_reg[230].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[230].genblk1.genblk1.latch.q ;
 wire \shift_reg[231].genblk1.genblk1.latch.clk ;
 wire \shift_reg[231].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[231].genblk1.genblk1.latch.q ;
 wire \shift_reg[232].genblk1.genblk1.latch.clk ;
 wire \shift_reg[232].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[232].genblk1.genblk1.latch.q ;
 wire \shift_reg[233].genblk1.genblk1.latch.clk ;
 wire \shift_reg[233].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[233].genblk1.genblk1.latch.q ;
 wire \shift_reg[234].genblk1.genblk1.latch.clk ;
 wire \shift_reg[234].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[234].genblk1.genblk1.latch.q ;
 wire \shift_reg[235].genblk1.genblk1.latch.clk ;
 wire \shift_reg[235].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[235].genblk1.genblk1.latch.q ;
 wire \shift_reg[236].genblk1.genblk1.latch.clk ;
 wire \shift_reg[236].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[236].genblk1.genblk1.latch.q ;
 wire \shift_reg[237].genblk1.genblk1.latch.clk ;
 wire \shift_reg[237].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[237].genblk1.genblk1.latch.q ;
 wire \shift_reg[238].genblk1.genblk1.latch.clk ;
 wire \shift_reg[238].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[238].genblk1.genblk1.latch.q ;
 wire \shift_reg[239].genblk1.genblk1.latch.clk ;
 wire \shift_reg[239].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[239].genblk1.genblk1.latch.q ;
 wire \shift_reg[23].genblk1.genblk1.latch.clk ;
 wire \shift_reg[23].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[23].genblk1.genblk1.latch.q ;
 wire \shift_reg[240].genblk1.genblk1.latch.clk ;
 wire \shift_reg[240].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[240].genblk1.genblk1.latch.q ;
 wire \shift_reg[241].genblk1.genblk1.latch.clk ;
 wire \shift_reg[241].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[241].genblk1.genblk1.latch.q ;
 wire \shift_reg[242].genblk1.genblk1.latch.clk ;
 wire \shift_reg[242].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[242].genblk1.genblk1.latch.q ;
 wire \shift_reg[243].genblk1.genblk1.latch.clk ;
 wire \shift_reg[243].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[243].genblk1.genblk1.latch.q ;
 wire \shift_reg[244].genblk1.genblk1.latch.clk ;
 wire \shift_reg[244].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[244].genblk1.genblk1.latch.q ;
 wire \shift_reg[245].genblk1.genblk1.latch.clk ;
 wire \shift_reg[245].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[245].genblk1.genblk1.latch.q ;
 wire \shift_reg[246].genblk1.genblk1.latch.clk ;
 wire \shift_reg[246].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[246].genblk1.genblk1.latch.q ;
 wire \shift_reg[247].genblk1.genblk1.latch.clk ;
 wire \shift_reg[247].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[247].genblk1.genblk1.latch.q ;
 wire \shift_reg[248].genblk1.genblk1.latch.clk ;
 wire \shift_reg[248].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[248].genblk1.genblk1.latch.q ;
 wire \shift_reg[249].genblk1.genblk1.latch.clk ;
 wire \shift_reg[249].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[249].genblk1.genblk1.latch.q ;
 wire \shift_reg[24].genblk1.genblk1.latch.clk ;
 wire \shift_reg[24].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[24].genblk1.genblk1.latch.q ;
 wire \shift_reg[250].genblk1.genblk1.latch.clk ;
 wire \shift_reg[250].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[250].genblk1.genblk1.latch.q ;
 wire \shift_reg[251].genblk1.genblk1.latch.clk ;
 wire \shift_reg[251].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[251].genblk1.genblk1.latch.q ;
 wire \shift_reg[252].genblk1.genblk1.latch.clk ;
 wire \shift_reg[252].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[252].genblk1.genblk1.latch.q ;
 wire \shift_reg[253].genblk1.genblk1.latch.clk ;
 wire \shift_reg[253].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[253].genblk1.genblk1.latch.q ;
 wire \shift_reg[254].genblk1.genblk1.latch.clk ;
 wire \shift_reg[254].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[254].genblk1.genblk1.latch.q ;
 wire \shift_reg[255].genblk1.genblk1.latch.clk ;
 wire \shift_reg[255].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[255].genblk1.genblk1.latch.q ;
 wire \shift_reg[256].genblk1.genblk1.latch.clk ;
 wire \shift_reg[256].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[256].genblk1.genblk1.latch.q ;
 wire \shift_reg[257].genblk1.genblk1.latch.clk ;
 wire \shift_reg[257].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[257].genblk1.genblk1.latch.q ;
 wire \shift_reg[258].genblk1.genblk1.latch.clk ;
 wire \shift_reg[258].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[258].genblk1.genblk1.latch.q ;
 wire \shift_reg[259].genblk1.genblk1.latch.clk ;
 wire \shift_reg[259].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[259].genblk1.genblk1.latch.q ;
 wire \shift_reg[25].genblk1.genblk1.latch.clk ;
 wire \shift_reg[25].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[25].genblk1.genblk1.latch.q ;
 wire \shift_reg[260].genblk1.genblk1.latch.clk ;
 wire \shift_reg[260].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[260].genblk1.genblk1.latch.q ;
 wire \shift_reg[261].genblk1.genblk1.latch.clk ;
 wire \shift_reg[261].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[261].genblk1.genblk1.latch.q ;
 wire \shift_reg[262].genblk1.genblk1.latch.clk ;
 wire \shift_reg[262].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[262].genblk1.genblk1.latch.q ;
 wire \shift_reg[263].genblk1.genblk1.latch.clk ;
 wire \shift_reg[263].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[263].genblk1.genblk1.latch.q ;
 wire \shift_reg[264].genblk1.genblk1.latch.clk ;
 wire \shift_reg[264].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[264].genblk1.genblk1.latch.q ;
 wire \shift_reg[265].genblk1.genblk1.latch.clk ;
 wire \shift_reg[265].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[265].genblk1.genblk1.latch.q ;
 wire \shift_reg[266].genblk1.genblk1.latch.clk ;
 wire \shift_reg[266].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[266].genblk1.genblk1.latch.q ;
 wire \shift_reg[267].genblk1.genblk1.latch.clk ;
 wire \shift_reg[267].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[267].genblk1.genblk1.latch.q ;
 wire \shift_reg[268].genblk1.genblk1.latch.clk ;
 wire \shift_reg[268].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[268].genblk1.genblk1.latch.q ;
 wire \shift_reg[269].genblk1.genblk1.latch.clk ;
 wire \shift_reg[269].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[269].genblk1.genblk1.latch.q ;
 wire \shift_reg[26].genblk1.genblk1.latch.clk ;
 wire \shift_reg[26].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[26].genblk1.genblk1.latch.q ;
 wire \shift_reg[270].genblk1.genblk1.latch.clk ;
 wire \shift_reg[270].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[270].genblk1.genblk1.latch.q ;
 wire \shift_reg[271].genblk1.genblk1.latch.clk ;
 wire \shift_reg[271].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[271].genblk1.genblk1.latch.q ;
 wire \shift_reg[272].genblk1.genblk1.latch.clk ;
 wire \shift_reg[272].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[272].genblk1.genblk1.latch.q ;
 wire \shift_reg[273].genblk1.genblk1.latch.clk ;
 wire \shift_reg[273].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[273].genblk1.genblk1.latch.q ;
 wire \shift_reg[274].genblk1.genblk1.latch.clk ;
 wire \shift_reg[274].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[274].genblk1.genblk1.latch.q ;
 wire \shift_reg[275].genblk1.genblk1.latch.clk ;
 wire \shift_reg[275].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[275].genblk1.genblk1.latch.q ;
 wire \shift_reg[276].genblk1.genblk1.latch.clk ;
 wire \shift_reg[276].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[276].genblk1.genblk1.latch.q ;
 wire \shift_reg[277].genblk1.genblk1.latch.clk ;
 wire \shift_reg[277].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[277].genblk1.genblk1.latch.q ;
 wire \shift_reg[278].genblk1.genblk1.latch.clk ;
 wire \shift_reg[278].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[278].genblk1.genblk1.latch.q ;
 wire \shift_reg[279].genblk1.genblk1.latch.clk ;
 wire \shift_reg[279].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[279].genblk1.genblk1.latch.q ;
 wire \shift_reg[27].genblk1.genblk1.latch.clk ;
 wire \shift_reg[27].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[27].genblk1.genblk1.latch.q ;
 wire \shift_reg[280].genblk1.genblk1.latch.clk ;
 wire \shift_reg[280].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[280].genblk1.genblk1.latch.q ;
 wire \shift_reg[281].genblk1.genblk1.latch.clk ;
 wire \shift_reg[281].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[281].genblk1.genblk1.latch.q ;
 wire \shift_reg[282].genblk1.genblk1.latch.clk ;
 wire \shift_reg[282].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[282].genblk1.genblk1.latch.q ;
 wire \shift_reg[283].genblk1.genblk1.latch.clk ;
 wire \shift_reg[283].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[283].genblk1.genblk1.latch.q ;
 wire \shift_reg[284].genblk1.genblk1.latch.clk ;
 wire \shift_reg[284].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[284].genblk1.genblk1.latch.q ;
 wire \shift_reg[285].genblk1.genblk1.latch.clk ;
 wire \shift_reg[285].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[285].genblk1.genblk1.latch.q ;
 wire \shift_reg[286].genblk1.genblk1.latch.clk ;
 wire \shift_reg[286].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[286].genblk1.genblk1.latch.q ;
 wire \shift_reg[287].genblk1.genblk1.latch.clk ;
 wire \shift_reg[287].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[287].genblk1.genblk1.latch.q ;
 wire \shift_reg[288].genblk1.genblk1.latch.clk ;
 wire \shift_reg[288].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[288].genblk1.genblk1.latch.q ;
 wire \shift_reg[289].genblk1.genblk1.latch.clk ;
 wire \shift_reg[289].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[289].genblk1.genblk1.latch.q ;
 wire \shift_reg[28].genblk1.genblk1.latch.clk ;
 wire \shift_reg[28].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[28].genblk1.genblk1.latch.q ;
 wire \shift_reg[290].genblk1.genblk1.latch.clk ;
 wire \shift_reg[290].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[290].genblk1.genblk1.latch.q ;
 wire \shift_reg[291].genblk1.genblk1.latch.clk ;
 wire \shift_reg[291].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[291].genblk1.genblk1.latch.q ;
 wire \shift_reg[292].genblk1.genblk1.latch.clk ;
 wire \shift_reg[292].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[292].genblk1.genblk1.latch.q ;
 wire \shift_reg[293].genblk1.genblk1.latch.clk ;
 wire \shift_reg[293].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[293].genblk1.genblk1.latch.q ;
 wire \shift_reg[294].genblk1.genblk1.latch.clk ;
 wire \shift_reg[294].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[294].genblk1.genblk1.latch.q ;
 wire \shift_reg[295].genblk1.genblk1.latch.clk ;
 wire \shift_reg[295].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[295].genblk1.genblk1.latch.q ;
 wire \shift_reg[296].genblk1.genblk1.latch.clk ;
 wire \shift_reg[296].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[296].genblk1.genblk1.latch.q ;
 wire \shift_reg[297].genblk1.genblk1.latch.clk ;
 wire \shift_reg[297].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[297].genblk1.genblk1.latch.q ;
 wire \shift_reg[298].genblk1.genblk1.latch.clk ;
 wire \shift_reg[298].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[298].genblk1.genblk1.latch.q ;
 wire \shift_reg[299].genblk1.genblk1.latch.clk ;
 wire \shift_reg[299].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[299].genblk1.genblk1.latch.q ;
 wire \shift_reg[29].genblk1.genblk1.latch.clk ;
 wire \shift_reg[29].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[29].genblk1.genblk1.latch.q ;
 wire \shift_reg[2].genblk1.genblk1.latch.clk ;
 wire \shift_reg[2].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[2].genblk1.genblk1.latch.q ;
 wire \shift_reg[300].genblk1.genblk1.latch.clk ;
 wire \shift_reg[300].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[300].genblk1.genblk1.latch.q ;
 wire \shift_reg[301].genblk1.genblk1.latch.clk ;
 wire \shift_reg[301].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[301].genblk1.genblk1.latch.q ;
 wire \shift_reg[302].genblk1.genblk1.latch.clk ;
 wire \shift_reg[302].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[302].genblk1.genblk1.latch.q ;
 wire \shift_reg[303].genblk1.genblk1.latch.clk ;
 wire \shift_reg[303].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[303].genblk1.genblk1.latch.q ;
 wire \shift_reg[304].genblk1.genblk1.latch.clk ;
 wire \shift_reg[304].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[304].genblk1.genblk1.latch.q ;
 wire \shift_reg[305].genblk1.genblk1.latch.clk ;
 wire \shift_reg[305].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[305].genblk1.genblk1.latch.q ;
 wire \shift_reg[306].genblk1.genblk1.latch.clk ;
 wire \shift_reg[306].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[306].genblk1.genblk1.latch.q ;
 wire \shift_reg[307].genblk1.genblk1.latch.clk ;
 wire \shift_reg[307].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[307].genblk1.genblk1.latch.q ;
 wire \shift_reg[308].genblk1.genblk1.latch.clk ;
 wire \shift_reg[308].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[308].genblk1.genblk1.latch.q ;
 wire \shift_reg[309].genblk1.genblk1.latch.clk ;
 wire \shift_reg[309].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[309].genblk1.genblk1.latch.q ;
 wire \shift_reg[30].genblk1.genblk1.latch.clk ;
 wire \shift_reg[30].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[30].genblk1.genblk1.latch.q ;
 wire \shift_reg[310].genblk1.genblk1.latch.clk ;
 wire \shift_reg[310].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[310].genblk1.genblk1.latch.q ;
 wire \shift_reg[311].genblk1.genblk1.latch.clk ;
 wire \shift_reg[311].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[311].genblk1.genblk1.latch.q ;
 wire \shift_reg[312].genblk1.genblk1.latch.clk ;
 wire \shift_reg[312].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[312].genblk1.genblk1.latch.q ;
 wire \shift_reg[313].genblk1.genblk1.latch.clk ;
 wire \shift_reg[313].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[313].genblk1.genblk1.latch.q ;
 wire \shift_reg[314].genblk1.genblk1.latch.clk ;
 wire \shift_reg[314].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[314].genblk1.genblk1.latch.q ;
 wire \shift_reg[315].genblk1.genblk1.latch.clk ;
 wire \shift_reg[315].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[315].genblk1.genblk1.latch.q ;
 wire \shift_reg[316].genblk1.genblk1.latch.clk ;
 wire \shift_reg[316].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[316].genblk1.genblk1.latch.q ;
 wire \shift_reg[317].genblk1.genblk1.latch.clk ;
 wire \shift_reg[317].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[317].genblk1.genblk1.latch.q ;
 wire \shift_reg[318].genblk1.genblk1.latch.clk ;
 wire \shift_reg[318].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[318].genblk1.genblk1.latch.q ;
 wire \shift_reg[319].genblk1.genblk1.latch.clk ;
 wire \shift_reg[319].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[319].genblk1.genblk1.latch.q ;
 wire \shift_reg[31].genblk1.genblk1.latch.clk ;
 wire \shift_reg[31].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[31].genblk1.genblk1.latch.q ;
 wire \shift_reg[320].genblk1.genblk1.latch.clk ;
 wire \shift_reg[320].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[320].genblk1.genblk1.latch.q ;
 wire \shift_reg[321].genblk1.genblk1.latch.clk ;
 wire \shift_reg[321].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[321].genblk1.genblk1.latch.q ;
 wire \shift_reg[322].genblk1.genblk1.latch.clk ;
 wire \shift_reg[322].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[322].genblk1.genblk1.latch.q ;
 wire \shift_reg[323].genblk1.genblk1.latch.clk ;
 wire \shift_reg[323].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[323].genblk1.genblk1.latch.q ;
 wire \shift_reg[324].genblk1.genblk1.latch.clk ;
 wire \shift_reg[324].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[324].genblk1.genblk1.latch.q ;
 wire \shift_reg[325].genblk1.genblk1.latch.clk ;
 wire \shift_reg[325].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[325].genblk1.genblk1.latch.q ;
 wire \shift_reg[326].genblk1.genblk1.latch.clk ;
 wire \shift_reg[326].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[326].genblk1.genblk1.latch.q ;
 wire \shift_reg[327].genblk1.genblk1.latch.clk ;
 wire \shift_reg[327].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[327].genblk1.genblk1.latch.q ;
 wire \shift_reg[328].genblk1.genblk1.latch.clk ;
 wire \shift_reg[328].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[328].genblk1.genblk1.latch.q ;
 wire \shift_reg[329].genblk1.genblk1.latch.clk ;
 wire \shift_reg[329].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[329].genblk1.genblk1.latch.q ;
 wire \shift_reg[32].genblk1.genblk1.latch.clk ;
 wire \shift_reg[32].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[32].genblk1.genblk1.latch.q ;
 wire \shift_reg[330].genblk1.genblk1.latch.clk ;
 wire \shift_reg[330].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[330].genblk1.genblk1.latch.q ;
 wire \shift_reg[331].genblk1.genblk1.latch.clk ;
 wire \shift_reg[331].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[331].genblk1.genblk1.latch.q ;
 wire \shift_reg[332].genblk1.genblk1.latch.clk ;
 wire \shift_reg[332].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[332].genblk1.genblk1.latch.q ;
 wire \shift_reg[333].genblk1.genblk1.latch.clk ;
 wire \shift_reg[333].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[333].genblk1.genblk1.latch.q ;
 wire \shift_reg[334].genblk1.genblk1.latch.clk ;
 wire \shift_reg[334].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[334].genblk1.genblk1.latch.q ;
 wire \shift_reg[335].genblk1.genblk1.latch.clk ;
 wire \shift_reg[335].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[335].genblk1.genblk1.latch.q ;
 wire \shift_reg[336].genblk1.genblk1.latch.clk ;
 wire \shift_reg[336].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[336].genblk1.genblk1.latch.q ;
 wire \shift_reg[337].genblk1.genblk1.latch.clk ;
 wire \shift_reg[337].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[337].genblk1.genblk1.latch.q ;
 wire \shift_reg[338].genblk1.genblk1.latch.clk ;
 wire \shift_reg[338].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[338].genblk1.genblk1.latch.q ;
 wire \shift_reg[339].genblk1.genblk1.latch.clk ;
 wire \shift_reg[339].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[339].genblk1.genblk1.latch.q ;
 wire \shift_reg[33].genblk1.genblk1.latch.clk ;
 wire \shift_reg[33].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[33].genblk1.genblk1.latch.q ;
 wire \shift_reg[340].genblk1.genblk1.latch.clk ;
 wire \shift_reg[340].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[340].genblk1.genblk1.latch.q ;
 wire \shift_reg[341].genblk1.genblk1.latch.clk ;
 wire \shift_reg[341].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[341].genblk1.genblk1.latch.q ;
 wire \shift_reg[342].genblk1.genblk1.latch.clk ;
 wire \shift_reg[342].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[342].genblk1.genblk1.latch.q ;
 wire \shift_reg[343].genblk1.genblk1.latch.clk ;
 wire \shift_reg[343].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[343].genblk1.genblk1.latch.q ;
 wire \shift_reg[344].genblk1.genblk1.latch.clk ;
 wire \shift_reg[344].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[344].genblk1.genblk1.latch.q ;
 wire \shift_reg[345].genblk1.genblk1.latch.clk ;
 wire \shift_reg[345].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[345].genblk1.genblk1.latch.q ;
 wire \shift_reg[346].genblk1.genblk1.latch.clk ;
 wire \shift_reg[346].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[346].genblk1.genblk1.latch.q ;
 wire \shift_reg[347].genblk1.genblk1.latch.clk ;
 wire \shift_reg[347].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[347].genblk1.genblk1.latch.q ;
 wire \shift_reg[348].genblk1.genblk1.latch.clk ;
 wire \shift_reg[348].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[348].genblk1.genblk1.latch.q ;
 wire \shift_reg[349].genblk1.genblk1.latch.clk ;
 wire \shift_reg[349].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[349].genblk1.genblk1.latch.q ;
 wire \shift_reg[34].genblk1.genblk1.latch.clk ;
 wire \shift_reg[34].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[34].genblk1.genblk1.latch.q ;
 wire \shift_reg[350].genblk1.genblk1.latch.clk ;
 wire \shift_reg[350].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[350].genblk1.genblk1.latch.q ;
 wire \shift_reg[351].genblk1.genblk1.latch.clk ;
 wire \shift_reg[351].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[351].genblk1.genblk1.latch.q ;
 wire \shift_reg[352].genblk1.genblk1.latch.clk ;
 wire \shift_reg[352].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[352].genblk1.genblk1.latch.q ;
 wire \shift_reg[353].genblk1.genblk1.latch.clk ;
 wire \shift_reg[353].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[353].genblk1.genblk1.latch.q ;
 wire \shift_reg[354].genblk1.genblk1.latch.clk ;
 wire \shift_reg[354].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[354].genblk1.genblk1.latch.q ;
 wire \shift_reg[355].genblk1.genblk1.latch.clk ;
 wire \shift_reg[355].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[355].genblk1.genblk1.latch.q ;
 wire \shift_reg[356].genblk1.genblk1.latch.clk ;
 wire \shift_reg[356].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[356].genblk1.genblk1.latch.q ;
 wire \shift_reg[357].genblk1.genblk1.latch.clk ;
 wire \shift_reg[357].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[357].genblk1.genblk1.latch.q ;
 wire \shift_reg[358].genblk1.genblk1.latch.clk ;
 wire \shift_reg[358].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[358].genblk1.genblk1.latch.q ;
 wire \shift_reg[359].genblk1.genblk1.latch.clk ;
 wire \shift_reg[359].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[359].genblk1.genblk1.latch.q ;
 wire \shift_reg[35].genblk1.genblk1.latch.clk ;
 wire \shift_reg[35].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[35].genblk1.genblk1.latch.q ;
 wire \shift_reg[360].genblk1.genblk1.latch.clk ;
 wire \shift_reg[360].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[360].genblk1.genblk1.latch.q ;
 wire \shift_reg[361].genblk1.genblk1.latch.clk ;
 wire \shift_reg[361].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[361].genblk1.genblk1.latch.q ;
 wire \shift_reg[362].genblk1.genblk1.latch.clk ;
 wire \shift_reg[362].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[362].genblk1.genblk1.latch.q ;
 wire \shift_reg[363].genblk1.genblk1.latch.clk ;
 wire \shift_reg[363].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[363].genblk1.genblk1.latch.q ;
 wire \shift_reg[364].genblk1.genblk1.latch.clk ;
 wire \shift_reg[364].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[364].genblk1.genblk1.latch.q ;
 wire \shift_reg[365].genblk1.genblk1.latch.clk ;
 wire \shift_reg[365].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[365].genblk1.genblk1.latch.q ;
 wire \shift_reg[366].genblk1.genblk1.latch.clk ;
 wire \shift_reg[366].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[366].genblk1.genblk1.latch.q ;
 wire \shift_reg[367].genblk1.genblk1.latch.clk ;
 wire \shift_reg[367].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[367].genblk1.genblk1.latch.q ;
 wire \shift_reg[368].genblk1.genblk1.latch.clk ;
 wire \shift_reg[368].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[368].genblk1.genblk1.latch.q ;
 wire \shift_reg[369].genblk1.genblk1.latch.clk ;
 wire \shift_reg[369].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[369].genblk1.genblk1.latch.q ;
 wire \shift_reg[36].genblk1.genblk1.latch.clk ;
 wire \shift_reg[36].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[36].genblk1.genblk1.latch.q ;
 wire \shift_reg[370].genblk1.genblk1.latch.clk ;
 wire \shift_reg[370].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[370].genblk1.genblk1.latch.q ;
 wire \shift_reg[371].genblk1.genblk1.latch.clk ;
 wire \shift_reg[371].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[371].genblk1.genblk1.latch.q ;
 wire \shift_reg[372].genblk1.genblk1.latch.clk ;
 wire \shift_reg[372].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[372].genblk1.genblk1.latch.q ;
 wire \shift_reg[373].genblk1.genblk1.latch.clk ;
 wire \shift_reg[373].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[373].genblk1.genblk1.latch.q ;
 wire \shift_reg[374].genblk1.genblk1.latch.clk ;
 wire \shift_reg[374].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[374].genblk1.genblk1.latch.q ;
 wire \shift_reg[375].genblk1.genblk1.latch.clk ;
 wire \shift_reg[375].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[375].genblk1.genblk1.latch.q ;
 wire \shift_reg[376].genblk1.genblk1.latch.clk ;
 wire \shift_reg[376].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[376].genblk1.genblk1.latch.q ;
 wire \shift_reg[377].genblk1.genblk1.latch.clk ;
 wire \shift_reg[377].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[377].genblk1.genblk1.latch.q ;
 wire \shift_reg[378].genblk1.genblk1.latch.clk ;
 wire \shift_reg[378].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[378].genblk1.genblk1.latch.q ;
 wire \shift_reg[379].genblk1.genblk1.latch.clk ;
 wire \shift_reg[379].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[379].genblk1.genblk1.latch.q ;
 wire \shift_reg[37].genblk1.genblk1.latch.clk ;
 wire \shift_reg[37].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[37].genblk1.genblk1.latch.q ;
 wire \shift_reg[380].genblk1.genblk1.latch.clk ;
 wire \shift_reg[380].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[380].genblk1.genblk1.latch.q ;
 wire \shift_reg[381].genblk1.genblk1.latch.clk ;
 wire \shift_reg[381].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[381].genblk1.genblk1.latch.q ;
 wire \shift_reg[382].genblk1.genblk1.latch.clk ;
 wire \shift_reg[382].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[382].genblk1.genblk1.latch.q ;
 wire \shift_reg[383].genblk1.genblk1.latch.clk ;
 wire \shift_reg[383].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[383].genblk1.genblk1.latch.q ;
 wire \shift_reg[384].genblk1.genblk1.latch.clk ;
 wire \shift_reg[384].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[384].genblk1.genblk1.latch.q ;
 wire \shift_reg[385].genblk1.genblk1.latch.clk ;
 wire \shift_reg[385].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[385].genblk1.genblk1.latch.q ;
 wire \shift_reg[386].genblk1.genblk1.latch.clk ;
 wire \shift_reg[386].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[386].genblk1.genblk1.latch.q ;
 wire \shift_reg[387].genblk1.genblk1.latch.clk ;
 wire \shift_reg[387].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[387].genblk1.genblk1.latch.q ;
 wire \shift_reg[388].genblk1.genblk1.latch.clk ;
 wire \shift_reg[388].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[388].genblk1.genblk1.latch.q ;
 wire \shift_reg[389].genblk1.genblk1.latch.clk ;
 wire \shift_reg[389].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[389].genblk1.genblk1.latch.q ;
 wire \shift_reg[38].genblk1.genblk1.latch.clk ;
 wire \shift_reg[38].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[38].genblk1.genblk1.latch.q ;
 wire \shift_reg[390].genblk1.genblk1.latch.clk ;
 wire \shift_reg[390].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[390].genblk1.genblk1.latch.q ;
 wire \shift_reg[391].genblk1.genblk1.latch.clk ;
 wire \shift_reg[391].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[391].genblk1.genblk1.latch.q ;
 wire \shift_reg[392].genblk1.genblk1.latch.clk ;
 wire \shift_reg[392].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[392].genblk1.genblk1.latch.q ;
 wire \shift_reg[393].genblk1.genblk1.latch.clk ;
 wire \shift_reg[393].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[393].genblk1.genblk1.latch.q ;
 wire \shift_reg[394].genblk1.genblk1.latch.clk ;
 wire \shift_reg[394].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[394].genblk1.genblk1.latch.q ;
 wire \shift_reg[395].genblk1.genblk1.latch.clk ;
 wire \shift_reg[395].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[395].genblk1.genblk1.latch.q ;
 wire \shift_reg[396].genblk1.genblk1.latch.clk ;
 wire \shift_reg[396].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[396].genblk1.genblk1.latch.q ;
 wire \shift_reg[397].genblk1.genblk1.latch.clk ;
 wire \shift_reg[397].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[397].genblk1.genblk1.latch.q ;
 wire \shift_reg[398].genblk1.genblk1.latch.clk ;
 wire \shift_reg[398].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[398].genblk1.genblk1.latch.q ;
 wire \shift_reg[399].genblk1.genblk1.latch.clk ;
 wire \shift_reg[399].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[399].genblk1.genblk1.latch.q ;
 wire \shift_reg[39].genblk1.genblk1.latch.clk ;
 wire \shift_reg[39].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[39].genblk1.genblk1.latch.q ;
 wire \shift_reg[3].genblk1.genblk1.latch.clk ;
 wire \shift_reg[3].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[3].genblk1.genblk1.latch.q ;
 wire \shift_reg[400].genblk1.genblk1.latch.clk ;
 wire \shift_reg[400].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[400].genblk1.genblk1.latch.q ;
 wire \shift_reg[401].genblk1.genblk1.latch.clk ;
 wire \shift_reg[401].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[401].genblk1.genblk1.latch.q ;
 wire \shift_reg[402].genblk1.genblk1.latch.clk ;
 wire \shift_reg[402].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[402].genblk1.genblk1.latch.q ;
 wire \shift_reg[403].genblk1.genblk1.latch.clk ;
 wire \shift_reg[403].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[403].genblk1.genblk1.latch.q ;
 wire \shift_reg[404].genblk1.genblk1.latch.clk ;
 wire \shift_reg[404].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[404].genblk1.genblk1.latch.q ;
 wire \shift_reg[405].genblk1.genblk1.latch.clk ;
 wire \shift_reg[405].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[405].genblk1.genblk1.latch.q ;
 wire \shift_reg[406].genblk1.genblk1.latch.clk ;
 wire \shift_reg[406].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[406].genblk1.genblk1.latch.q ;
 wire \shift_reg[407].genblk1.genblk1.latch.clk ;
 wire \shift_reg[407].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[407].genblk1.genblk1.latch.q ;
 wire \shift_reg[408].genblk1.genblk1.latch.clk ;
 wire \shift_reg[408].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[408].genblk1.genblk1.latch.q ;
 wire \shift_reg[409].genblk1.genblk1.latch.clk ;
 wire \shift_reg[409].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[409].genblk1.genblk1.latch.q ;
 wire \shift_reg[40].genblk1.genblk1.latch.clk ;
 wire \shift_reg[40].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[40].genblk1.genblk1.latch.q ;
 wire \shift_reg[410].genblk1.genblk1.latch.clk ;
 wire \shift_reg[410].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[410].genblk1.genblk1.latch.q ;
 wire \shift_reg[411].genblk1.genblk1.latch.clk ;
 wire \shift_reg[411].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[411].genblk1.genblk1.latch.q ;
 wire \shift_reg[412].genblk1.genblk1.latch.clk ;
 wire \shift_reg[412].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[412].genblk1.genblk1.latch.q ;
 wire \shift_reg[413].genblk1.genblk1.latch.clk ;
 wire \shift_reg[413].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[413].genblk1.genblk1.latch.q ;
 wire \shift_reg[414].genblk1.genblk1.latch.clk ;
 wire \shift_reg[414].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[414].genblk1.genblk1.latch.q ;
 wire \shift_reg[415].genblk1.genblk1.latch.clk ;
 wire \shift_reg[415].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[415].genblk1.genblk1.latch.q ;
 wire \shift_reg[416].genblk1.genblk1.latch.clk ;
 wire \shift_reg[416].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[416].genblk1.genblk1.latch.q ;
 wire \shift_reg[417].genblk1.genblk1.latch.clk ;
 wire \shift_reg[417].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[417].genblk1.genblk1.latch.q ;
 wire \shift_reg[418].genblk1.genblk1.latch.clk ;
 wire \shift_reg[418].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[418].genblk1.genblk1.latch.q ;
 wire \shift_reg[419].genblk1.genblk1.latch.clk ;
 wire \shift_reg[419].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[419].genblk1.genblk1.latch.q ;
 wire \shift_reg[41].genblk1.genblk1.latch.clk ;
 wire \shift_reg[41].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[41].genblk1.genblk1.latch.q ;
 wire \shift_reg[420].genblk1.genblk1.latch.clk ;
 wire \shift_reg[420].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[420].genblk1.genblk1.latch.q ;
 wire \shift_reg[421].genblk1.genblk1.latch.clk ;
 wire \shift_reg[421].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[421].genblk1.genblk1.latch.q ;
 wire \shift_reg[422].genblk1.genblk1.latch.clk ;
 wire \shift_reg[422].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[422].genblk1.genblk1.latch.q ;
 wire \shift_reg[423].genblk1.genblk1.latch.clk ;
 wire \shift_reg[423].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[423].genblk1.genblk1.latch.q ;
 wire \shift_reg[424].genblk1.genblk1.latch.clk ;
 wire \shift_reg[424].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[424].genblk1.genblk1.latch.q ;
 wire \shift_reg[425].genblk1.genblk1.latch.clk ;
 wire \shift_reg[425].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[425].genblk1.genblk1.latch.q ;
 wire \shift_reg[426].genblk1.genblk1.latch.clk ;
 wire \shift_reg[426].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[426].genblk1.genblk1.latch.q ;
 wire \shift_reg[427].genblk1.genblk1.latch.clk ;
 wire \shift_reg[427].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[427].genblk1.genblk1.latch.q ;
 wire \shift_reg[428].genblk1.genblk1.latch.clk ;
 wire \shift_reg[428].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[428].genblk1.genblk1.latch.q ;
 wire \shift_reg[429].genblk1.genblk1.latch.clk ;
 wire \shift_reg[429].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[429].genblk1.genblk1.latch.q ;
 wire \shift_reg[42].genblk1.genblk1.latch.clk ;
 wire \shift_reg[42].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[42].genblk1.genblk1.latch.q ;
 wire \shift_reg[430].genblk1.genblk1.latch.clk ;
 wire \shift_reg[430].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[430].genblk1.genblk1.latch.q ;
 wire \shift_reg[431].genblk1.genblk1.latch.clk ;
 wire \shift_reg[431].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[431].genblk1.genblk1.latch.q ;
 wire \shift_reg[432].genblk1.genblk1.latch.clk ;
 wire \shift_reg[432].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[432].genblk1.genblk1.latch.q ;
 wire \shift_reg[433].genblk1.genblk1.latch.clk ;
 wire \shift_reg[433].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[433].genblk1.genblk1.latch.q ;
 wire \shift_reg[434].genblk1.genblk1.latch.clk ;
 wire \shift_reg[434].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[434].genblk1.genblk1.latch.q ;
 wire \shift_reg[435].genblk1.genblk1.latch.clk ;
 wire \shift_reg[435].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[435].genblk1.genblk1.latch.q ;
 wire \shift_reg[436].genblk1.genblk1.latch.clk ;
 wire \shift_reg[436].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[436].genblk1.genblk1.latch.q ;
 wire \shift_reg[437].genblk1.genblk1.latch.clk ;
 wire \shift_reg[437].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[437].genblk1.genblk1.latch.q ;
 wire \shift_reg[438].genblk1.genblk1.latch.clk ;
 wire \shift_reg[438].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[438].genblk1.genblk1.latch.q ;
 wire \shift_reg[439].genblk1.genblk1.latch.clk ;
 wire \shift_reg[439].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[439].genblk1.genblk1.latch.q ;
 wire \shift_reg[43].genblk1.genblk1.latch.clk ;
 wire \shift_reg[43].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[43].genblk1.genblk1.latch.q ;
 wire \shift_reg[440].genblk1.genblk1.latch.clk ;
 wire \shift_reg[440].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[440].genblk1.genblk1.latch.q ;
 wire \shift_reg[441].genblk1.genblk1.latch.clk ;
 wire \shift_reg[441].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[441].genblk1.genblk1.latch.q ;
 wire \shift_reg[442].genblk1.genblk1.latch.clk ;
 wire \shift_reg[442].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[442].genblk1.genblk1.latch.q ;
 wire \shift_reg[443].genblk1.genblk1.latch.clk ;
 wire \shift_reg[443].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[443].genblk1.genblk1.latch.q ;
 wire \shift_reg[444].genblk1.genblk1.latch.clk ;
 wire \shift_reg[444].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[444].genblk1.genblk1.latch.q ;
 wire \shift_reg[445].genblk1.genblk1.latch.clk ;
 wire \shift_reg[445].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[445].genblk1.genblk1.latch.q ;
 wire \shift_reg[446].genblk1.genblk1.latch.clk ;
 wire \shift_reg[446].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[446].genblk1.genblk1.latch.q ;
 wire \shift_reg[447].genblk1.genblk1.latch.clk ;
 wire \shift_reg[447].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[447].genblk1.genblk1.latch.q ;
 wire \shift_reg[448].genblk1.genblk1.latch.clk ;
 wire \shift_reg[448].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[448].genblk1.genblk1.latch.q ;
 wire \shift_reg[449].genblk1.genblk1.latch.clk ;
 wire \shift_reg[449].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[449].genblk1.genblk1.latch.q ;
 wire \shift_reg[44].genblk1.genblk1.latch.clk ;
 wire \shift_reg[44].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[44].genblk1.genblk1.latch.q ;
 wire \shift_reg[450].genblk1.genblk1.latch.clk ;
 wire \shift_reg[450].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[450].genblk1.genblk1.latch.q ;
 wire \shift_reg[451].genblk1.genblk1.latch.clk ;
 wire \shift_reg[451].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[451].genblk1.genblk1.latch.q ;
 wire \shift_reg[452].genblk1.genblk1.latch.clk ;
 wire \shift_reg[452].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[452].genblk1.genblk1.latch.q ;
 wire \shift_reg[453].genblk1.genblk1.latch.clk ;
 wire \shift_reg[453].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[453].genblk1.genblk1.latch.q ;
 wire \shift_reg[454].genblk1.genblk1.latch.clk ;
 wire \shift_reg[454].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[454].genblk1.genblk1.latch.q ;
 wire \shift_reg[455].genblk1.genblk1.latch.clk ;
 wire \shift_reg[455].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[455].genblk1.genblk1.latch.q ;
 wire \shift_reg[456].genblk1.genblk1.latch.clk ;
 wire \shift_reg[456].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[456].genblk1.genblk1.latch.q ;
 wire \shift_reg[457].genblk1.genblk1.latch.clk ;
 wire \shift_reg[457].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[457].genblk1.genblk1.latch.q ;
 wire \shift_reg[458].genblk1.genblk1.latch.clk ;
 wire \shift_reg[458].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[458].genblk1.genblk1.latch.q ;
 wire \shift_reg[459].genblk1.genblk1.latch.clk ;
 wire \shift_reg[459].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[459].genblk1.genblk1.latch.q ;
 wire \shift_reg[45].genblk1.genblk1.latch.clk ;
 wire \shift_reg[45].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[45].genblk1.genblk1.latch.q ;
 wire \shift_reg[460].genblk1.genblk1.latch.clk ;
 wire \shift_reg[460].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[460].genblk1.genblk1.latch.q ;
 wire \shift_reg[461].genblk1.genblk1.latch.clk ;
 wire \shift_reg[461].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[461].genblk1.genblk1.latch.q ;
 wire \shift_reg[462].genblk1.genblk1.latch.clk ;
 wire \shift_reg[462].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[462].genblk1.genblk1.latch.q ;
 wire \shift_reg[463].genblk1.genblk1.latch.clk ;
 wire \shift_reg[463].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[463].genblk1.genblk1.latch.q ;
 wire \shift_reg[464].genblk1.genblk1.latch.clk ;
 wire \shift_reg[464].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[464].genblk1.genblk1.latch.q ;
 wire \shift_reg[465].genblk1.genblk1.latch.clk ;
 wire \shift_reg[465].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[465].genblk1.genblk1.latch.q ;
 wire \shift_reg[466].genblk1.genblk1.latch.clk ;
 wire \shift_reg[466].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[466].genblk1.genblk1.latch.q ;
 wire \shift_reg[467].genblk1.genblk1.latch.clk ;
 wire \shift_reg[467].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[467].genblk1.genblk1.latch.q ;
 wire \shift_reg[468].genblk1.genblk1.latch.clk ;
 wire \shift_reg[468].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[468].genblk1.genblk1.latch.q ;
 wire \shift_reg[469].genblk1.genblk1.latch.clk ;
 wire \shift_reg[469].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[469].genblk1.genblk1.latch.q ;
 wire \shift_reg[46].genblk1.genblk1.latch.clk ;
 wire \shift_reg[46].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[46].genblk1.genblk1.latch.q ;
 wire \shift_reg[470].genblk1.genblk1.latch.clk ;
 wire \shift_reg[470].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[470].genblk1.genblk1.latch.q ;
 wire \shift_reg[471].genblk1.genblk1.latch.clk ;
 wire \shift_reg[471].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[471].genblk1.genblk1.latch.q ;
 wire \shift_reg[472].genblk1.genblk1.latch.clk ;
 wire \shift_reg[472].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[472].genblk1.genblk1.latch.q ;
 wire \shift_reg[473].genblk1.genblk1.latch.clk ;
 wire \shift_reg[473].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[473].genblk1.genblk1.latch.q ;
 wire \shift_reg[474].genblk1.genblk1.latch.clk ;
 wire \shift_reg[474].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[474].genblk1.genblk1.latch.q ;
 wire \shift_reg[475].genblk1.genblk1.latch.clk ;
 wire \shift_reg[475].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[475].genblk1.genblk1.latch.q ;
 wire \shift_reg[476].genblk1.genblk1.latch.clk ;
 wire \shift_reg[476].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[476].genblk1.genblk1.latch.q ;
 wire \shift_reg[477].genblk1.genblk1.latch.clk ;
 wire \shift_reg[477].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[477].genblk1.genblk1.latch.q ;
 wire \shift_reg[478].genblk1.genblk1.latch.clk ;
 wire \shift_reg[478].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[478].genblk1.genblk1.latch.q ;
 wire \shift_reg[479].genblk1.genblk1.latch.clk ;
 wire \shift_reg[479].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[479].genblk1.genblk1.latch.q ;
 wire \shift_reg[47].genblk1.genblk1.latch.clk ;
 wire \shift_reg[47].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[47].genblk1.genblk1.latch.q ;
 wire \shift_reg[480].genblk1.genblk1.latch.clk ;
 wire \shift_reg[480].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[480].genblk1.genblk1.latch.q ;
 wire \shift_reg[481].genblk1.genblk1.latch.clk ;
 wire \shift_reg[481].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[481].genblk1.genblk1.latch.q ;
 wire \shift_reg[482].genblk1.genblk1.latch.clk ;
 wire \shift_reg[482].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[482].genblk1.genblk1.latch.q ;
 wire \shift_reg[483].genblk1.genblk1.latch.clk ;
 wire \shift_reg[483].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[483].genblk1.genblk1.latch.q ;
 wire \shift_reg[484].genblk1.genblk1.latch.clk ;
 wire \shift_reg[484].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[484].genblk1.genblk1.latch.q ;
 wire \shift_reg[485].genblk1.genblk1.latch.clk ;
 wire \shift_reg[485].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[485].genblk1.genblk1.latch.q ;
 wire \shift_reg[486].genblk1.genblk1.latch.clk ;
 wire \shift_reg[486].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[486].genblk1.genblk1.latch.q ;
 wire \shift_reg[487].genblk1.genblk1.latch.clk ;
 wire \shift_reg[487].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[487].genblk1.genblk1.latch.q ;
 wire \shift_reg[488].genblk1.genblk1.latch.clk ;
 wire \shift_reg[488].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[488].genblk1.genblk1.latch.q ;
 wire \shift_reg[489].genblk1.genblk1.latch.clk ;
 wire \shift_reg[489].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[489].genblk1.genblk1.latch.q ;
 wire \shift_reg[48].genblk1.genblk1.latch.clk ;
 wire \shift_reg[48].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[48].genblk1.genblk1.latch.q ;
 wire \shift_reg[490].genblk1.genblk1.latch.clk ;
 wire \shift_reg[490].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[490].genblk1.genblk1.latch.q ;
 wire \shift_reg[491].genblk1.genblk1.latch.clk ;
 wire \shift_reg[491].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[491].genblk1.genblk1.latch.q ;
 wire \shift_reg[492].genblk1.genblk1.latch.clk ;
 wire \shift_reg[492].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[492].genblk1.genblk1.latch.q ;
 wire \shift_reg[493].genblk1.genblk1.latch.clk ;
 wire \shift_reg[493].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[493].genblk1.genblk1.latch.q ;
 wire \shift_reg[494].genblk1.genblk1.latch.clk ;
 wire \shift_reg[494].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[494].genblk1.genblk1.latch.q ;
 wire \shift_reg[495].genblk1.genblk1.latch.clk ;
 wire \shift_reg[495].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[495].genblk1.genblk1.latch.q ;
 wire \shift_reg[496].genblk1.genblk1.latch.clk ;
 wire \shift_reg[496].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[496].genblk1.genblk1.latch.q ;
 wire \shift_reg[497].genblk1.genblk1.latch.clk ;
 wire \shift_reg[497].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[497].genblk1.genblk1.latch.q ;
 wire \shift_reg[498].genblk1.genblk1.latch.clk ;
 wire \shift_reg[498].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[498].genblk1.genblk1.latch.q ;
 wire \shift_reg[499].genblk1.genblk1.latch.clk ;
 wire \shift_reg[499].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[499].genblk1.genblk1.latch.q ;
 wire \shift_reg[49].genblk1.genblk1.latch.clk ;
 wire \shift_reg[49].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[49].genblk1.genblk1.latch.q ;
 wire \shift_reg[4].genblk1.genblk1.latch.clk ;
 wire \shift_reg[4].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[4].genblk1.genblk1.latch.q ;
 wire \shift_reg[500].genblk1.genblk1.latch.clk ;
 wire \shift_reg[500].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[500].genblk1.genblk1.latch.q ;
 wire \shift_reg[501].genblk1.genblk1.latch.clk ;
 wire \shift_reg[501].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[501].genblk1.genblk1.latch.q ;
 wire \shift_reg[502].genblk1.genblk1.latch.clk ;
 wire \shift_reg[502].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[502].genblk1.genblk1.latch.q ;
 wire \shift_reg[503].genblk1.genblk1.latch.clk ;
 wire \shift_reg[503].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[503].genblk1.genblk1.latch.q ;
 wire \shift_reg[504].genblk1.genblk1.latch.clk ;
 wire \shift_reg[504].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[504].genblk1.genblk1.latch.q ;
 wire \shift_reg[505].genblk1.genblk1.latch.clk ;
 wire \shift_reg[505].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[505].genblk1.genblk1.latch.q ;
 wire \shift_reg[506].genblk1.genblk1.latch.clk ;
 wire \shift_reg[506].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[506].genblk1.genblk1.latch.q ;
 wire \shift_reg[507].genblk1.genblk1.latch.clk ;
 wire \shift_reg[507].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[507].genblk1.genblk1.latch.q ;
 wire \shift_reg[508].genblk1.genblk1.latch.clk ;
 wire \shift_reg[508].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[508].genblk1.genblk1.latch.q ;
 wire \shift_reg[509].genblk1.genblk1.latch.clk ;
 wire \shift_reg[509].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[509].genblk1.genblk1.latch.q ;
 wire \shift_reg[50].genblk1.genblk1.latch.clk ;
 wire \shift_reg[50].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[50].genblk1.genblk1.latch.q ;
 wire \shift_reg[510].genblk1.genblk1.latch.clk ;
 wire \shift_reg[510].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[510].genblk1.genblk1.latch.q ;
 wire \shift_reg[511].genblk1.genblk1.latch.clk ;
 wire \shift_reg[511].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[511].genblk1.genblk1.latch.q ;
 wire \shift_reg[51].genblk1.genblk1.latch.clk ;
 wire \shift_reg[51].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[51].genblk1.genblk1.latch.q ;
 wire \shift_reg[52].genblk1.genblk1.latch.clk ;
 wire \shift_reg[52].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[52].genblk1.genblk1.latch.q ;
 wire \shift_reg[53].genblk1.genblk1.latch.clk ;
 wire \shift_reg[53].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[53].genblk1.genblk1.latch.q ;
 wire \shift_reg[54].genblk1.genblk1.latch.clk ;
 wire \shift_reg[54].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[54].genblk1.genblk1.latch.q ;
 wire \shift_reg[55].genblk1.genblk1.latch.clk ;
 wire \shift_reg[55].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[55].genblk1.genblk1.latch.q ;
 wire \shift_reg[56].genblk1.genblk1.latch.clk ;
 wire \shift_reg[56].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[56].genblk1.genblk1.latch.q ;
 wire \shift_reg[57].genblk1.genblk1.latch.clk ;
 wire \shift_reg[57].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[57].genblk1.genblk1.latch.q ;
 wire \shift_reg[58].genblk1.genblk1.latch.clk ;
 wire \shift_reg[58].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[58].genblk1.genblk1.latch.q ;
 wire \shift_reg[59].genblk1.genblk1.latch.clk ;
 wire \shift_reg[59].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[59].genblk1.genblk1.latch.q ;
 wire \shift_reg[5].genblk1.genblk1.latch.clk ;
 wire \shift_reg[5].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[5].genblk1.genblk1.latch.q ;
 wire \shift_reg[60].genblk1.genblk1.latch.clk ;
 wire \shift_reg[60].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[60].genblk1.genblk1.latch.q ;
 wire \shift_reg[61].genblk1.genblk1.latch.clk ;
 wire \shift_reg[61].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[61].genblk1.genblk1.latch.q ;
 wire \shift_reg[62].genblk1.genblk1.latch.clk ;
 wire \shift_reg[62].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[62].genblk1.genblk1.latch.q ;
 wire \shift_reg[63].genblk1.genblk1.latch.clk ;
 wire \shift_reg[63].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[63].genblk1.genblk1.latch.q ;
 wire \shift_reg[64].genblk1.genblk1.latch.clk ;
 wire \shift_reg[64].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[64].genblk1.genblk1.latch.q ;
 wire \shift_reg[65].genblk1.genblk1.latch.clk ;
 wire \shift_reg[65].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[65].genblk1.genblk1.latch.q ;
 wire \shift_reg[66].genblk1.genblk1.latch.clk ;
 wire \shift_reg[66].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[66].genblk1.genblk1.latch.q ;
 wire \shift_reg[67].genblk1.genblk1.latch.clk ;
 wire \shift_reg[67].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[67].genblk1.genblk1.latch.q ;
 wire \shift_reg[68].genblk1.genblk1.latch.clk ;
 wire \shift_reg[68].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[68].genblk1.genblk1.latch.q ;
 wire \shift_reg[69].genblk1.genblk1.latch.clk ;
 wire \shift_reg[69].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[69].genblk1.genblk1.latch.q ;
 wire \shift_reg[6].genblk1.genblk1.latch.clk ;
 wire \shift_reg[6].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[6].genblk1.genblk1.latch.q ;
 wire \shift_reg[70].genblk1.genblk1.latch.clk ;
 wire \shift_reg[70].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[70].genblk1.genblk1.latch.q ;
 wire \shift_reg[71].genblk1.genblk1.latch.clk ;
 wire \shift_reg[71].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[71].genblk1.genblk1.latch.q ;
 wire \shift_reg[72].genblk1.genblk1.latch.clk ;
 wire \shift_reg[72].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[72].genblk1.genblk1.latch.q ;
 wire \shift_reg[73].genblk1.genblk1.latch.clk ;
 wire \shift_reg[73].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[73].genblk1.genblk1.latch.q ;
 wire \shift_reg[74].genblk1.genblk1.latch.clk ;
 wire \shift_reg[74].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[74].genblk1.genblk1.latch.q ;
 wire \shift_reg[75].genblk1.genblk1.latch.clk ;
 wire \shift_reg[75].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[75].genblk1.genblk1.latch.q ;
 wire \shift_reg[76].genblk1.genblk1.latch.clk ;
 wire \shift_reg[76].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[76].genblk1.genblk1.latch.q ;
 wire \shift_reg[77].genblk1.genblk1.latch.clk ;
 wire \shift_reg[77].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[77].genblk1.genblk1.latch.q ;
 wire \shift_reg[78].genblk1.genblk1.latch.clk ;
 wire \shift_reg[78].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[78].genblk1.genblk1.latch.q ;
 wire \shift_reg[79].genblk1.genblk1.latch.clk ;
 wire \shift_reg[79].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[79].genblk1.genblk1.latch.q ;
 wire \shift_reg[7].genblk1.genblk1.latch.clk ;
 wire \shift_reg[7].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[7].genblk1.genblk1.latch.q ;
 wire \shift_reg[80].genblk1.genblk1.latch.clk ;
 wire \shift_reg[80].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[80].genblk1.genblk1.latch.q ;
 wire \shift_reg[81].genblk1.genblk1.latch.clk ;
 wire \shift_reg[81].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[81].genblk1.genblk1.latch.q ;
 wire \shift_reg[82].genblk1.genblk1.latch.clk ;
 wire \shift_reg[82].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[82].genblk1.genblk1.latch.q ;
 wire \shift_reg[83].genblk1.genblk1.latch.clk ;
 wire \shift_reg[83].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[83].genblk1.genblk1.latch.q ;
 wire \shift_reg[84].genblk1.genblk1.latch.clk ;
 wire \shift_reg[84].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[84].genblk1.genblk1.latch.q ;
 wire \shift_reg[85].genblk1.genblk1.latch.clk ;
 wire \shift_reg[85].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[85].genblk1.genblk1.latch.q ;
 wire \shift_reg[86].genblk1.genblk1.latch.clk ;
 wire \shift_reg[86].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[86].genblk1.genblk1.latch.q ;
 wire \shift_reg[87].genblk1.genblk1.latch.clk ;
 wire \shift_reg[87].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[87].genblk1.genblk1.latch.q ;
 wire \shift_reg[88].genblk1.genblk1.latch.clk ;
 wire \shift_reg[88].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[88].genblk1.genblk1.latch.q ;
 wire \shift_reg[89].genblk1.genblk1.latch.clk ;
 wire \shift_reg[89].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[89].genblk1.genblk1.latch.q ;
 wire \shift_reg[8].genblk1.genblk1.latch.clk ;
 wire \shift_reg[8].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[8].genblk1.genblk1.latch.q ;
 wire \shift_reg[90].genblk1.genblk1.latch.clk ;
 wire \shift_reg[90].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[90].genblk1.genblk1.latch.q ;
 wire \shift_reg[91].genblk1.genblk1.latch.clk ;
 wire \shift_reg[91].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[91].genblk1.genblk1.latch.q ;
 wire \shift_reg[92].genblk1.genblk1.latch.clk ;
 wire \shift_reg[92].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[92].genblk1.genblk1.latch.q ;
 wire \shift_reg[93].genblk1.genblk1.latch.clk ;
 wire \shift_reg[93].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[93].genblk1.genblk1.latch.q ;
 wire \shift_reg[94].genblk1.genblk1.latch.clk ;
 wire \shift_reg[94].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[94].genblk1.genblk1.latch.q ;
 wire \shift_reg[95].genblk1.genblk1.latch.clk ;
 wire \shift_reg[95].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[95].genblk1.genblk1.latch.q ;
 wire \shift_reg[96].genblk1.genblk1.latch.clk ;
 wire \shift_reg[96].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[96].genblk1.genblk1.latch.q ;
 wire \shift_reg[97].genblk1.genblk1.latch.clk ;
 wire \shift_reg[97].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[97].genblk1.genblk1.latch.q ;
 wire \shift_reg[98].genblk1.genblk1.latch.clk ;
 wire \shift_reg[98].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[98].genblk1.genblk1.latch.q ;
 wire \shift_reg[99].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[9].genblk1.genblk1.latch.nclk ;
 wire \u_invA.out ;
 wire \u_invB.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;

 sky130_fd_sc_hd__xor2_1 _000_ (.A(\u_invB.out ),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\shift_reg[511].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__dlxtp_1 _001_ (.D(\shift_reg[2].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[3].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[3].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _002_ (.D(\shift_reg[3].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[4].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[4].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _003_ (.D(\shift_reg[4].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[5].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[5].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _004_ (.D(\shift_reg[5].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[6].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[6].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _005_ (.D(\shift_reg[6].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[7].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[7].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _006_ (.D(\shift_reg[7].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[8].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[8].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _007_ (.D(\shift_reg[8].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[10].genblk1.genblk1.latch.clkout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[10].genblk1.genblk1.latch.d ));
 sky130_fd_sc_hd__dlxtp_1 _008_ (.D(\shift_reg[10].genblk1.genblk1.latch.d ),
    .GATE(\shift_reg[10].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[10].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _009_ (.D(\shift_reg[10].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[11].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[11].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _010_ (.D(\shift_reg[11].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[12].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[12].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _011_ (.D(\shift_reg[12].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[13].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[13].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _012_ (.D(\shift_reg[13].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[14].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[14].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _013_ (.D(\shift_reg[14].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[15].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[15].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _014_ (.D(\shift_reg[15].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[16].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[16].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _015_ (.D(\shift_reg[16].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[17].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[17].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _016_ (.D(\shift_reg[17].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[18].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[18].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _017_ (.D(\shift_reg[18].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[19].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[19].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _018_ (.D(\shift_reg[19].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[20].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[20].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _019_ (.D(\shift_reg[20].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[21].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[21].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _020_ (.D(\shift_reg[21].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[22].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[22].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _021_ (.D(\shift_reg[22].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[23].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[23].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _022_ (.D(\shift_reg[23].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[24].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[24].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _023_ (.D(\shift_reg[24].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[25].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[25].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _024_ (.D(\shift_reg[25].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[26].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[26].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _025_ (.D(\shift_reg[26].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[27].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[27].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _026_ (.D(\shift_reg[27].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[28].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[28].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _027_ (.D(\shift_reg[28].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[29].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[29].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _028_ (.D(\shift_reg[29].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[30].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[30].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _029_ (.D(\shift_reg[30].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[31].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[31].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _030_ (.D(\shift_reg[31].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[32].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[32].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _031_ (.D(\shift_reg[32].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[33].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[33].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _032_ (.D(\shift_reg[33].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[34].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[34].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _033_ (.D(\shift_reg[34].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[35].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[35].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _034_ (.D(\shift_reg[35].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[36].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[36].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _035_ (.D(\shift_reg[36].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[37].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[37].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _036_ (.D(\shift_reg[37].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[38].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[38].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _037_ (.D(\shift_reg[38].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[39].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[39].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _038_ (.D(\shift_reg[39].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[40].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[40].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _039_ (.D(\shift_reg[40].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[41].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[41].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _040_ (.D(\shift_reg[41].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[42].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[42].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _041_ (.D(\shift_reg[42].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[43].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[43].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _042_ (.D(\shift_reg[43].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[44].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[44].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _043_ (.D(\shift_reg[44].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[45].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[45].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _044_ (.D(\shift_reg[45].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[46].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[46].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _045_ (.D(\shift_reg[46].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[47].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[47].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _046_ (.D(\shift_reg[47].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[48].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[48].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _047_ (.D(\shift_reg[48].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[49].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[49].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _048_ (.D(\shift_reg[49].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[50].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[50].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _049_ (.D(\shift_reg[50].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[51].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[51].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _050_ (.D(\shift_reg[51].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[52].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[52].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _051_ (.D(\shift_reg[52].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[53].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[53].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _052_ (.D(\shift_reg[53].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[54].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[54].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _053_ (.D(\shift_reg[54].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[55].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[55].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _054_ (.D(\shift_reg[55].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[56].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[56].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _055_ (.D(\shift_reg[56].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[57].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[57].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _056_ (.D(\shift_reg[57].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[58].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[58].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _057_ (.D(\shift_reg[58].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[59].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[59].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _058_ (.D(\shift_reg[59].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[60].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[60].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _059_ (.D(\shift_reg[60].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[61].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[61].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _060_ (.D(\shift_reg[61].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[62].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[62].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _061_ (.D(\shift_reg[62].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[63].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[63].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _062_ (.D(\shift_reg[63].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[64].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[64].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _063_ (.D(\shift_reg[64].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[65].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[65].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _064_ (.D(\shift_reg[65].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[66].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[66].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _065_ (.D(\shift_reg[66].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[67].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[67].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _066_ (.D(\shift_reg[67].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[68].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[68].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _067_ (.D(\shift_reg[68].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[69].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[69].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _068_ (.D(\shift_reg[69].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[70].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[70].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _069_ (.D(\shift_reg[70].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[71].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[71].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _070_ (.D(\shift_reg[71].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[72].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[72].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _071_ (.D(\shift_reg[72].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[73].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[73].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _072_ (.D(\shift_reg[73].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[74].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[74].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _073_ (.D(\shift_reg[74].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[75].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[75].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _074_ (.D(\shift_reg[75].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[76].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[76].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _075_ (.D(\shift_reg[76].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[77].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[77].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _076_ (.D(\shift_reg[77].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[78].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[78].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _077_ (.D(\shift_reg[78].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[79].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[79].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _078_ (.D(\shift_reg[79].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[80].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[80].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _079_ (.D(\shift_reg[80].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[81].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[81].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _080_ (.D(\shift_reg[81].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[82].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[82].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _081_ (.D(\shift_reg[82].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[83].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[83].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _082_ (.D(\shift_reg[83].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[84].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[84].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _083_ (.D(\shift_reg[84].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[85].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[85].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _084_ (.D(\shift_reg[85].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[86].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[86].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _085_ (.D(\shift_reg[86].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[87].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[87].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _086_ (.D(\shift_reg[87].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[88].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[88].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _087_ (.D(\shift_reg[88].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[89].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[89].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _088_ (.D(\shift_reg[89].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[90].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[90].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _089_ (.D(\shift_reg[90].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[91].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[91].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _090_ (.D(\shift_reg[91].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[92].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[92].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _091_ (.D(\shift_reg[92].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[93].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[93].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _092_ (.D(\shift_reg[93].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[94].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[94].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _093_ (.D(\shift_reg[94].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[95].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[95].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _094_ (.D(\shift_reg[95].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[96].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[96].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _095_ (.D(\shift_reg[96].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[97].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[97].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _096_ (.D(\shift_reg[97].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[98].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[98].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _097_ (.D(\shift_reg[98].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[100].genblk1.genblk1.latch.clkout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[100].genblk1.genblk1.latch.d ));
 sky130_fd_sc_hd__dlxtp_1 _098_ (.D(\shift_reg[100].genblk1.genblk1.latch.d ),
    .GATE(\shift_reg[100].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[100].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _099_ (.D(\shift_reg[100].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[101].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[101].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _100_ (.D(\shift_reg[101].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[102].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[102].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _101_ (.D(\shift_reg[102].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[103].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[103].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _102_ (.D(\shift_reg[103].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[104].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[104].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _103_ (.D(\shift_reg[104].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[105].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[105].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _104_ (.D(\shift_reg[105].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[106].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[106].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _105_ (.D(\shift_reg[106].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[107].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[107].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _106_ (.D(\shift_reg[107].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[108].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[108].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _107_ (.D(\shift_reg[108].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[109].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[109].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _108_ (.D(\shift_reg[109].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[110].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[110].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _109_ (.D(\shift_reg[110].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[111].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[111].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _110_ (.D(\shift_reg[111].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[112].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[112].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _111_ (.D(\shift_reg[112].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[113].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[113].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _112_ (.D(\shift_reg[113].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[114].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[114].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _113_ (.D(\shift_reg[114].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[115].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[115].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _114_ (.D(\shift_reg[115].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[116].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[116].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _115_ (.D(\shift_reg[116].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[117].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[117].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _116_ (.D(\shift_reg[117].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[118].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[118].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _117_ (.D(\shift_reg[118].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[119].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[119].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _118_ (.D(\shift_reg[119].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[120].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[120].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _119_ (.D(\shift_reg[120].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[121].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[121].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _120_ (.D(\shift_reg[121].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[122].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[122].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _121_ (.D(\shift_reg[122].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[123].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[123].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _122_ (.D(\shift_reg[123].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[124].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[124].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _123_ (.D(\shift_reg[124].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[125].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[125].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _124_ (.D(\shift_reg[125].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[126].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[126].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _125_ (.D(\shift_reg[126].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[127].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[127].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _126_ (.D(\shift_reg[127].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[128].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[128].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _127_ (.D(\shift_reg[128].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[129].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[129].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _128_ (.D(\shift_reg[129].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[130].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[130].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _129_ (.D(\shift_reg[130].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[131].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[131].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _130_ (.D(\shift_reg[131].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[132].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[132].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _131_ (.D(\shift_reg[132].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[133].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[133].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _132_ (.D(\shift_reg[133].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[134].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[134].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _133_ (.D(\shift_reg[134].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[135].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[135].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _134_ (.D(\shift_reg[135].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[136].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[136].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _135_ (.D(\shift_reg[136].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[137].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[137].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _136_ (.D(\shift_reg[137].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[138].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[138].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _137_ (.D(\shift_reg[138].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[139].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[139].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _138_ (.D(\shift_reg[139].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[140].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[140].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _139_ (.D(\shift_reg[140].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[141].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[141].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _140_ (.D(\shift_reg[141].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[142].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[142].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _141_ (.D(\shift_reg[142].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[143].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[143].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _142_ (.D(\shift_reg[143].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[144].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[144].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _143_ (.D(\shift_reg[144].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[145].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[145].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _144_ (.D(\shift_reg[145].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[146].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[146].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _145_ (.D(\shift_reg[146].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[147].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[147].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _146_ (.D(\shift_reg[147].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[148].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[148].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _147_ (.D(\shift_reg[148].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[149].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[149].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _148_ (.D(\shift_reg[149].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[150].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[150].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _149_ (.D(\shift_reg[150].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[151].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[151].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _150_ (.D(\shift_reg[151].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[152].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[152].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _151_ (.D(\shift_reg[152].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[153].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[153].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _152_ (.D(\shift_reg[153].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[154].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[154].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _153_ (.D(\shift_reg[154].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[155].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[155].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _154_ (.D(\shift_reg[155].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[156].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[156].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _155_ (.D(\shift_reg[156].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[157].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[157].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _156_ (.D(\shift_reg[157].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[158].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[158].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _157_ (.D(\shift_reg[158].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[159].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[159].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _158_ (.D(\shift_reg[159].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[160].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[160].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _159_ (.D(\shift_reg[160].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[161].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[161].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _160_ (.D(\shift_reg[161].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[162].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[162].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _161_ (.D(\shift_reg[162].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[163].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[163].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _162_ (.D(\shift_reg[163].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[164].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[164].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _163_ (.D(\shift_reg[164].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[165].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[165].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _164_ (.D(\shift_reg[165].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[166].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[166].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _165_ (.D(\shift_reg[166].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[167].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[167].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _166_ (.D(\shift_reg[167].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[168].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[168].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _167_ (.D(\shift_reg[168].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[169].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[169].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _168_ (.D(\shift_reg[169].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[170].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[170].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _169_ (.D(\shift_reg[170].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[171].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[171].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _170_ (.D(\shift_reg[171].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[172].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[172].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _171_ (.D(\shift_reg[172].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[173].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[173].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _172_ (.D(\shift_reg[173].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[174].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[174].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _173_ (.D(\shift_reg[174].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[175].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[175].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _174_ (.D(\shift_reg[175].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[176].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[176].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _175_ (.D(\shift_reg[176].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[177].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[177].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _176_ (.D(\shift_reg[177].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[178].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[178].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _177_ (.D(\shift_reg[178].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[179].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[179].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _178_ (.D(\shift_reg[179].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[180].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[180].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _179_ (.D(\shift_reg[180].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[181].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[181].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _180_ (.D(\shift_reg[181].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[182].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[182].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _181_ (.D(\shift_reg[182].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[183].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[183].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _182_ (.D(\shift_reg[183].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[184].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[184].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _183_ (.D(\shift_reg[184].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[185].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[185].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _184_ (.D(\shift_reg[185].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[186].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[186].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _185_ (.D(\shift_reg[186].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[187].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[187].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _186_ (.D(\shift_reg[187].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[188].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[188].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _187_ (.D(\shift_reg[188].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[189].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[189].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _188_ (.D(\shift_reg[189].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[190].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[190].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _189_ (.D(\shift_reg[190].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[191].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[191].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _190_ (.D(\shift_reg[191].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[192].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[192].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _191_ (.D(\shift_reg[192].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[193].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[193].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _192_ (.D(\shift_reg[193].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[194].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[194].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _193_ (.D(\shift_reg[194].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[195].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[195].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _194_ (.D(\shift_reg[195].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[196].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[196].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _195_ (.D(\shift_reg[196].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[197].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[197].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _196_ (.D(\shift_reg[197].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[198].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[198].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _197_ (.D(\shift_reg[198].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[199].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[199].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _198_ (.D(\shift_reg[199].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[200].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[200].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _199_ (.D(\shift_reg[200].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[201].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[201].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _200_ (.D(\shift_reg[201].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[202].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[202].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _201_ (.D(\shift_reg[202].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[203].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[203].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _202_ (.D(\shift_reg[203].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[204].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[204].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _203_ (.D(\shift_reg[204].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[205].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[205].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _204_ (.D(\shift_reg[205].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[206].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[206].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _205_ (.D(\shift_reg[206].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[207].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[207].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _206_ (.D(\shift_reg[207].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[208].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[208].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _207_ (.D(\shift_reg[208].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[209].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[209].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _208_ (.D(\shift_reg[209].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[210].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[210].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _209_ (.D(\shift_reg[210].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[211].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[211].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _210_ (.D(\shift_reg[211].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[212].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[212].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _211_ (.D(\shift_reg[212].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[213].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[213].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _212_ (.D(\shift_reg[213].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[214].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[214].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _213_ (.D(\shift_reg[214].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[215].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[215].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _214_ (.D(\shift_reg[215].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[216].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[216].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _215_ (.D(\shift_reg[216].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[217].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[217].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _216_ (.D(\shift_reg[217].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[218].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[218].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _217_ (.D(\shift_reg[218].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[219].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[219].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _218_ (.D(\shift_reg[219].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[220].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[220].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _219_ (.D(\shift_reg[220].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[221].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[221].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _220_ (.D(\shift_reg[221].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[222].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[222].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _221_ (.D(\shift_reg[222].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[223].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[223].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _222_ (.D(\shift_reg[223].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[224].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[224].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _223_ (.D(\shift_reg[224].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[225].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[225].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _224_ (.D(\shift_reg[225].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[226].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[226].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _225_ (.D(\shift_reg[226].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[227].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[227].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _226_ (.D(\shift_reg[227].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[228].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[228].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _227_ (.D(\shift_reg[228].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[229].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[229].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _228_ (.D(\shift_reg[229].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[230].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[230].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _229_ (.D(\shift_reg[230].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[231].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[231].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _230_ (.D(\shift_reg[231].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[232].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[232].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _231_ (.D(\shift_reg[232].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[233].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[233].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _232_ (.D(\shift_reg[233].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[234].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[234].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _233_ (.D(\shift_reg[234].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[235].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[235].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _234_ (.D(\shift_reg[235].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[236].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[236].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _235_ (.D(\shift_reg[236].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[237].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[237].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _236_ (.D(\shift_reg[237].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[238].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[238].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _237_ (.D(\shift_reg[238].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[239].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[239].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _238_ (.D(\shift_reg[239].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[240].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[240].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _239_ (.D(\shift_reg[240].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[241].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[241].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _240_ (.D(\shift_reg[241].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[242].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[242].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _241_ (.D(\shift_reg[242].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[243].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[243].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _242_ (.D(\shift_reg[243].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[244].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[244].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _243_ (.D(\shift_reg[244].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[245].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[245].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _244_ (.D(\shift_reg[245].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[246].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[246].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _245_ (.D(\shift_reg[246].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[247].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[247].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _246_ (.D(\shift_reg[247].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[248].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[248].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _247_ (.D(\shift_reg[248].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[249].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[249].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _248_ (.D(\shift_reg[249].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[250].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[250].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _249_ (.D(\shift_reg[250].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[251].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[251].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _250_ (.D(\shift_reg[251].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[252].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[252].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _251_ (.D(\shift_reg[252].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[253].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[253].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _252_ (.D(\shift_reg[253].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[254].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[254].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _253_ (.D(\shift_reg[254].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[255].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[255].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _254_ (.D(\shift_reg[255].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[256].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[256].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _255_ (.D(\shift_reg[256].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[257].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[257].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _256_ (.D(\shift_reg[257].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[258].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[258].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _257_ (.D(\shift_reg[258].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[259].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[259].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _258_ (.D(\shift_reg[259].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[260].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[260].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _259_ (.D(\shift_reg[260].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[261].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[261].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _260_ (.D(\shift_reg[261].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[262].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[262].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _261_ (.D(\shift_reg[262].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[263].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[263].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _262_ (.D(\shift_reg[263].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[264].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[264].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _263_ (.D(\shift_reg[264].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[265].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[265].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _264_ (.D(\shift_reg[265].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[266].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[266].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _265_ (.D(\shift_reg[266].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[267].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[267].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _266_ (.D(\shift_reg[267].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[268].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[268].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _267_ (.D(\shift_reg[268].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[269].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[269].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _268_ (.D(\shift_reg[269].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[270].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[270].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _269_ (.D(\shift_reg[270].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[271].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[271].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _270_ (.D(\shift_reg[271].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[272].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[272].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _271_ (.D(\shift_reg[272].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[273].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[273].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _272_ (.D(\shift_reg[273].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[274].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[274].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _273_ (.D(\shift_reg[274].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[275].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[275].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _274_ (.D(\shift_reg[275].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[276].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[276].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _275_ (.D(\shift_reg[276].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[277].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[277].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _276_ (.D(\shift_reg[277].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[278].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[278].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _277_ (.D(\shift_reg[278].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[279].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[279].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _278_ (.D(\shift_reg[279].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[280].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[280].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _279_ (.D(\shift_reg[280].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[281].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[281].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _280_ (.D(\shift_reg[281].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[282].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[282].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _281_ (.D(\shift_reg[282].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[283].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[283].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _282_ (.D(\shift_reg[283].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[284].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[284].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _283_ (.D(\shift_reg[284].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[285].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[285].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _284_ (.D(\shift_reg[285].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[286].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[286].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _285_ (.D(\shift_reg[286].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[287].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[287].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _286_ (.D(\shift_reg[287].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[288].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[288].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _287_ (.D(\shift_reg[288].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[289].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[289].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _288_ (.D(\shift_reg[289].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[290].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[290].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _289_ (.D(\shift_reg[290].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[291].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[291].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _290_ (.D(\shift_reg[291].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[292].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[292].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _291_ (.D(\shift_reg[292].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[293].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[293].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _292_ (.D(\shift_reg[293].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[294].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[294].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _293_ (.D(\shift_reg[294].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[295].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[295].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _294_ (.D(\shift_reg[295].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[296].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[296].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _295_ (.D(\shift_reg[296].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[297].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[297].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _296_ (.D(\shift_reg[297].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[298].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[298].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _297_ (.D(\shift_reg[298].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[299].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[299].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _298_ (.D(\shift_reg[299].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[300].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[300].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _299_ (.D(\shift_reg[300].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[301].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[301].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _300_ (.D(\shift_reg[301].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[302].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[302].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _301_ (.D(\shift_reg[302].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[303].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[303].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _302_ (.D(\shift_reg[303].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[304].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[304].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _303_ (.D(\shift_reg[304].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[305].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[305].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _304_ (.D(\shift_reg[305].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[306].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[306].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _305_ (.D(\shift_reg[306].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[307].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[307].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _306_ (.D(\shift_reg[307].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[308].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[308].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _307_ (.D(\shift_reg[308].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[309].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[309].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _308_ (.D(\shift_reg[309].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[310].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[310].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _309_ (.D(\shift_reg[310].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[311].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[311].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _310_ (.D(\shift_reg[311].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[312].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[312].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _311_ (.D(\shift_reg[312].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[313].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[313].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _312_ (.D(\shift_reg[313].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[314].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[314].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _313_ (.D(\shift_reg[314].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[315].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[315].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _314_ (.D(\shift_reg[315].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[316].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[316].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _315_ (.D(\shift_reg[316].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[317].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[317].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _316_ (.D(\shift_reg[317].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[318].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[318].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _317_ (.D(\shift_reg[318].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[319].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[319].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _318_ (.D(\shift_reg[319].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[320].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[320].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _319_ (.D(\shift_reg[320].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[321].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[321].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _320_ (.D(\shift_reg[321].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[322].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[322].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _321_ (.D(\shift_reg[322].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[323].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[323].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _322_ (.D(\shift_reg[323].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[324].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[324].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _323_ (.D(\shift_reg[324].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[325].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[325].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _324_ (.D(\shift_reg[325].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[326].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[326].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _325_ (.D(\shift_reg[326].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[327].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[327].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _326_ (.D(\shift_reg[327].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[328].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[328].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _327_ (.D(\shift_reg[328].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[329].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[329].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _328_ (.D(\shift_reg[329].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[330].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[330].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _329_ (.D(\shift_reg[330].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[331].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[331].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _330_ (.D(\shift_reg[331].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[332].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[332].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _331_ (.D(\shift_reg[332].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[333].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[333].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _332_ (.D(\shift_reg[333].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[334].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[334].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _333_ (.D(\shift_reg[334].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[335].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[335].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _334_ (.D(\shift_reg[335].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[336].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[336].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _335_ (.D(\shift_reg[336].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[337].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[337].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _336_ (.D(\shift_reg[337].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[338].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[338].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _337_ (.D(\shift_reg[338].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[339].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[339].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _338_ (.D(\shift_reg[339].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[340].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[340].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _339_ (.D(\shift_reg[340].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[341].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[341].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _340_ (.D(\shift_reg[341].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[342].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[342].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _341_ (.D(\shift_reg[342].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[343].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[343].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _342_ (.D(\shift_reg[343].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[344].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[344].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _343_ (.D(\shift_reg[344].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[345].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[345].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _344_ (.D(\shift_reg[345].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[346].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[346].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _345_ (.D(\shift_reg[346].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[347].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[347].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _346_ (.D(\shift_reg[347].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[348].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[348].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _347_ (.D(\shift_reg[348].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[349].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[349].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _348_ (.D(\shift_reg[349].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[350].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[350].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _349_ (.D(\shift_reg[350].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[351].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[351].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _350_ (.D(\shift_reg[351].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[352].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[352].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _351_ (.D(\shift_reg[352].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[353].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[353].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _352_ (.D(\shift_reg[353].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[354].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[354].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _353_ (.D(\shift_reg[354].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[355].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[355].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _354_ (.D(\shift_reg[355].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[356].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[356].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _355_ (.D(\shift_reg[356].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[357].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[357].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _356_ (.D(\shift_reg[357].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[358].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[358].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _357_ (.D(\shift_reg[358].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[359].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[359].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _358_ (.D(\shift_reg[359].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[360].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[360].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _359_ (.D(\shift_reg[360].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[361].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[361].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _360_ (.D(\shift_reg[361].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[362].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[362].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _361_ (.D(\shift_reg[362].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[363].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[363].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _362_ (.D(\shift_reg[363].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[364].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[364].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _363_ (.D(\shift_reg[364].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[365].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[365].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _364_ (.D(\shift_reg[365].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[366].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[366].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _365_ (.D(\shift_reg[366].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[367].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[367].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _366_ (.D(\shift_reg[367].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[368].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[368].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _367_ (.D(\shift_reg[368].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[369].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[369].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _368_ (.D(\shift_reg[369].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[370].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[370].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _369_ (.D(\shift_reg[370].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[371].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[371].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _370_ (.D(\shift_reg[371].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[372].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[372].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _371_ (.D(\shift_reg[372].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[373].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[373].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _372_ (.D(\shift_reg[373].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[374].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[374].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _373_ (.D(\shift_reg[374].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[375].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[375].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _374_ (.D(\shift_reg[375].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[376].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[376].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _375_ (.D(\shift_reg[376].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[377].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[377].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _376_ (.D(\shift_reg[377].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[378].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[378].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _377_ (.D(\shift_reg[378].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[379].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[379].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _378_ (.D(\shift_reg[379].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[380].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[380].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _379_ (.D(\shift_reg[380].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[381].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[381].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _380_ (.D(\shift_reg[381].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[382].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[382].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _381_ (.D(\shift_reg[382].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[383].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[383].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _382_ (.D(\shift_reg[383].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[384].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[384].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _383_ (.D(\shift_reg[384].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[385].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[385].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _384_ (.D(\shift_reg[385].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[386].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[386].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _385_ (.D(\shift_reg[386].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[387].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[387].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _386_ (.D(\shift_reg[387].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[388].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[388].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _387_ (.D(\shift_reg[388].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[389].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[389].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _388_ (.D(\shift_reg[389].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[390].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[390].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _389_ (.D(\shift_reg[390].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[391].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[391].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _390_ (.D(\shift_reg[391].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[392].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[392].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _391_ (.D(\shift_reg[392].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[393].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[393].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _392_ (.D(\shift_reg[393].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[394].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[394].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _393_ (.D(\shift_reg[394].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[395].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[395].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _394_ (.D(\shift_reg[395].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[396].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[396].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _395_ (.D(\shift_reg[396].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[397].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[397].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _396_ (.D(\shift_reg[397].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[398].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[398].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _397_ (.D(\shift_reg[398].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[399].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[399].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _398_ (.D(\shift_reg[399].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[400].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[400].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _399_ (.D(\shift_reg[400].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[401].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[401].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _400_ (.D(\shift_reg[401].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[402].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[402].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _401_ (.D(\shift_reg[402].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[403].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[403].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _402_ (.D(\shift_reg[403].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[404].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[404].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _403_ (.D(\shift_reg[404].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[405].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[405].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _404_ (.D(\shift_reg[405].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[406].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[406].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _405_ (.D(\shift_reg[406].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[407].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[407].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _406_ (.D(\shift_reg[407].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[408].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[408].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _407_ (.D(\shift_reg[408].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[409].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[409].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _408_ (.D(\shift_reg[409].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[410].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[410].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _409_ (.D(\shift_reg[410].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[411].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[411].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _410_ (.D(\shift_reg[411].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[412].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[412].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _411_ (.D(\shift_reg[412].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[413].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[413].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _412_ (.D(\shift_reg[413].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[414].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[414].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _413_ (.D(\shift_reg[414].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[415].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[415].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _414_ (.D(\shift_reg[415].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[416].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[416].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _415_ (.D(\shift_reg[416].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[417].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[417].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _416_ (.D(\shift_reg[417].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[418].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[418].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _417_ (.D(\shift_reg[418].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[419].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[419].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _418_ (.D(\shift_reg[419].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[420].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[420].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _419_ (.D(\shift_reg[420].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[421].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[421].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _420_ (.D(\shift_reg[421].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[422].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[422].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _421_ (.D(\shift_reg[422].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[423].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[423].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _422_ (.D(\shift_reg[423].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[424].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[424].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _423_ (.D(\shift_reg[424].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[425].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[425].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _424_ (.D(\shift_reg[425].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[426].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[426].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _425_ (.D(\shift_reg[426].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[427].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[427].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _426_ (.D(\shift_reg[427].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[428].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[428].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _427_ (.D(\shift_reg[428].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[429].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[429].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _428_ (.D(\shift_reg[429].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[430].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[430].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _429_ (.D(\shift_reg[430].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[431].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[431].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _430_ (.D(\shift_reg[431].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[432].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[432].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _431_ (.D(\shift_reg[432].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[433].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[433].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _432_ (.D(\shift_reg[433].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[434].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[434].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _433_ (.D(\shift_reg[434].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[435].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[435].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _434_ (.D(\shift_reg[435].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[436].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[436].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _435_ (.D(\shift_reg[436].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[437].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[437].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _436_ (.D(\shift_reg[437].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[438].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[438].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _437_ (.D(\shift_reg[438].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[439].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[439].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _438_ (.D(\shift_reg[439].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[440].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[440].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _439_ (.D(\shift_reg[440].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[441].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[441].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _440_ (.D(\shift_reg[441].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[442].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[442].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _441_ (.D(\shift_reg[442].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[443].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[443].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _442_ (.D(\shift_reg[443].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[444].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[444].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _443_ (.D(\shift_reg[444].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[445].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[445].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _444_ (.D(\shift_reg[445].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[446].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[446].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _445_ (.D(\shift_reg[446].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[447].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[447].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _446_ (.D(\shift_reg[447].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[448].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[448].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _447_ (.D(\shift_reg[448].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[449].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[449].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _448_ (.D(\shift_reg[449].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[450].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[450].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _449_ (.D(\shift_reg[450].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[451].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[451].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _450_ (.D(\shift_reg[451].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[452].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[452].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _451_ (.D(\shift_reg[452].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[453].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[453].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _452_ (.D(\shift_reg[453].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[454].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[454].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _453_ (.D(\shift_reg[454].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[455].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[455].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _454_ (.D(\shift_reg[455].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[456].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[456].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _455_ (.D(\shift_reg[456].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[457].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[457].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _456_ (.D(\shift_reg[457].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[458].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[458].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _457_ (.D(\shift_reg[458].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[459].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[459].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _458_ (.D(\shift_reg[459].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[460].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[460].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _459_ (.D(\shift_reg[460].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[461].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[461].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _460_ (.D(\shift_reg[461].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[462].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[462].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _461_ (.D(\shift_reg[462].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[463].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[463].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _462_ (.D(\shift_reg[463].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[464].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[464].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _463_ (.D(\shift_reg[464].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[465].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[465].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _464_ (.D(\shift_reg[465].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[466].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[466].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _465_ (.D(\shift_reg[466].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[467].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[467].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _466_ (.D(\shift_reg[467].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[468].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[468].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _467_ (.D(\shift_reg[468].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[469].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[469].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _468_ (.D(\shift_reg[469].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[470].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[470].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _469_ (.D(\shift_reg[470].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[471].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[471].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _470_ (.D(\shift_reg[471].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[472].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[472].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _471_ (.D(\shift_reg[472].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[473].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[473].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _472_ (.D(\shift_reg[473].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[474].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[474].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _473_ (.D(\shift_reg[474].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[475].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[475].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _474_ (.D(\shift_reg[475].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[476].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[476].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _475_ (.D(\shift_reg[476].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[477].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[477].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _476_ (.D(\shift_reg[477].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[478].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[478].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _477_ (.D(\shift_reg[478].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[479].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[479].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _478_ (.D(\shift_reg[479].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[480].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[480].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _479_ (.D(\shift_reg[480].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[481].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[481].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _480_ (.D(\shift_reg[481].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[482].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[482].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _481_ (.D(\shift_reg[482].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[483].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[483].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _482_ (.D(\shift_reg[483].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[484].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[484].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _483_ (.D(\shift_reg[484].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[485].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[485].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _484_ (.D(\shift_reg[485].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[486].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[486].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _485_ (.D(\shift_reg[486].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[487].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[487].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _486_ (.D(\shift_reg[487].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[488].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[488].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _487_ (.D(\shift_reg[488].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[489].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[489].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _488_ (.D(\shift_reg[489].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[490].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[490].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _489_ (.D(\shift_reg[490].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[491].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[491].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _490_ (.D(\shift_reg[491].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[492].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[492].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _491_ (.D(\shift_reg[492].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[493].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[493].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _492_ (.D(\shift_reg[493].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[494].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[494].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _493_ (.D(\shift_reg[494].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[495].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[495].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _494_ (.D(\shift_reg[495].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[496].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[496].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _495_ (.D(\shift_reg[496].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[497].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[497].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _496_ (.D(\shift_reg[497].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[498].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[498].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _497_ (.D(\shift_reg[498].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[499].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[499].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _498_ (.D(\shift_reg[499].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[500].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[500].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _499_ (.D(\shift_reg[500].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[501].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[501].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _500_ (.D(\shift_reg[501].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[502].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[502].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _501_ (.D(\shift_reg[502].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[503].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[503].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _502_ (.D(\shift_reg[503].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[504].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[504].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _503_ (.D(\shift_reg[504].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[505].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[505].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _504_ (.D(\shift_reg[505].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[506].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[506].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _505_ (.D(\shift_reg[506].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[507].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[507].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _506_ (.D(\shift_reg[507].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[508].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[508].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _507_ (.D(\shift_reg[508].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[509].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[509].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _508_ (.D(\shift_reg[509].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[510].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[510].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _509_ (.D(\shift_reg[510].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[511].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[511].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _510_ (.D(net1),
    .GATE(\shift_reg[0].genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[0].genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _511_ (.D(\shift_reg[0].genblk1.latch.q ),
    .GATE(\shift_reg[1].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[1].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__dlxtp_1 _512_ (.D(\shift_reg[1].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[2].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_reg[2].genblk1.genblk1.latch.q ));
 sky130_fd_sc_hd__buf_2 _513_ (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _514_ (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _515_ (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _516_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__buf_2 _517_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__buf_2 _518_ (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__buf_2 _519_ (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _520_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__buf_2 _521_ (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__buf_2 _522_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _523_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__buf_2 _524_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__buf_2 _525_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__buf_2 _526_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__buf_2 _527_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _528_ (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__clkbuf_4 _529_ (.A(\shift_reg[511].genblk1.genblk1.latch.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _530_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _531_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _532_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _533_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _534_ (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _535_ (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _536_ (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_1 \shift_reg[100].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[100].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[100].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[100].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[100].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[100].genblk1.genblk1.latch.clkout ));
 sky130_fd_sc_hd__inv_1 \shift_reg[101].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[101].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[101].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[101].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[101].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[100].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[102].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[102].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[102].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[102].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[102].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[101].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[103].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[103].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[103].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[103].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[103].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[102].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[104].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[104].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[104].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[104].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[104].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[103].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[105].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[105].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[105].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[105].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[105].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[104].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[106].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[106].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[106].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[106].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[106].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[105].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[107].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[107].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[107].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[107].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[107].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[106].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[108].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[108].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[108].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[108].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[108].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[107].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[109].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[109].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[109].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[109].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[109].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[108].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[10].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[10].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[10].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[10].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[10].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[10].genblk1.genblk1.latch.clkout ));
 sky130_fd_sc_hd__inv_1 \shift_reg[110].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[110].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[110].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[110].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[110].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[109].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[111].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[111].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[111].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[111].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[111].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[110].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[112].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[112].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[112].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[112].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[112].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[111].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[113].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[113].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[113].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[113].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[113].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[112].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[114].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[114].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[114].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[114].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[114].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[113].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[115].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[115].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[115].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[115].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[115].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[114].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[116].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[116].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[116].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[116].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[116].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[115].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[117].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[117].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[117].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[117].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[117].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[116].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[118].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[118].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[118].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[118].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[118].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[117].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[119].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[119].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[119].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[119].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[119].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[118].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[11].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[11].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[11].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[11].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[11].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[10].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[120].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[120].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[120].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[120].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[120].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[119].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[121].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[121].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[121].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[121].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[121].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[120].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[122].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[122].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[122].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[122].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[122].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[121].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[123].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[123].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[123].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[123].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[123].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[122].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[124].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[124].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[124].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[124].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[124].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[123].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[125].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[125].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[125].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[125].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[125].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[124].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[126].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[126].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[126].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[126].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[126].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[125].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[127].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[127].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[127].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[127].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[127].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[126].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[128].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[128].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[128].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[128].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[128].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[127].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[129].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[129].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[129].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[129].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[129].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[128].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[12].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[12].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[12].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[12].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[12].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[11].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[130].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[130].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[130].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[130].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[130].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[129].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[131].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[131].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[131].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[131].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[131].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[130].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[132].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[132].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[132].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[132].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[132].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[131].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[133].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[133].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[133].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[133].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[133].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[132].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[134].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[134].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[134].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[134].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[134].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[133].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[135].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[135].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[135].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[135].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[135].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[134].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[136].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[136].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[136].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[136].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[136].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[135].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[137].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[137].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[137].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[137].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[137].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[136].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[138].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[138].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[138].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[138].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[138].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[137].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[139].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[139].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[139].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[139].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[139].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[138].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[13].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[13].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[13].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[13].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[13].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[12].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[140].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[140].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[140].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[140].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[140].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[139].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[141].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[141].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[141].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[141].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[141].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[140].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[142].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[142].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[142].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[142].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[142].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[141].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[143].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[143].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[143].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[143].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[143].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[142].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[144].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[144].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[144].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[144].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[144].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[143].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[145].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[145].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[145].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[145].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[145].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[144].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[146].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[146].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[146].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[146].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[146].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[145].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[147].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[147].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[147].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[147].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[147].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[146].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[148].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[148].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[148].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[148].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[148].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[147].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[149].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[149].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[149].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[149].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[149].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[148].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[14].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[14].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[14].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[14].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[14].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[13].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[150].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[150].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[150].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[150].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[150].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[149].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[151].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[151].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[151].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[151].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[151].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[150].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[152].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[152].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[152].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[152].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[152].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[151].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[153].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[153].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[153].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[153].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[153].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[152].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[154].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[154].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[154].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[154].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[154].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[153].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[155].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[155].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[155].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[155].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[155].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[154].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[156].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[156].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[156].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[156].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[156].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[155].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[157].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[157].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[157].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[157].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[157].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[156].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[158].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[158].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[158].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[158].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[158].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[157].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[159].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[159].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[159].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[159].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[159].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[158].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[15].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[15].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[15].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[15].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[15].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[14].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[160].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[160].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[160].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[160].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[160].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[159].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[161].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[161].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[161].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[161].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[161].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[160].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[162].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[162].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[162].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[162].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[162].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[161].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[163].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[163].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[163].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[163].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[163].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[162].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[164].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[164].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[164].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[164].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[164].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[163].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[165].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[165].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[165].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[165].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[165].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[164].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[166].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[166].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[166].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[166].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[166].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[165].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[167].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[167].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[167].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[167].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[167].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[166].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[168].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[168].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[168].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[168].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[168].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[167].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[169].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[169].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[169].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[169].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[169].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[168].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[16].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[16].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[16].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[16].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[16].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[15].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[170].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[170].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[170].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[170].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[170].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[169].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[171].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[171].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[171].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[171].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[171].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[170].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[172].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[172].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[172].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[172].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[172].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[171].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[173].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[173].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[173].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[173].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[173].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[172].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[174].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[174].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[174].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[174].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[174].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[173].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[175].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[175].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[175].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[175].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[175].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[174].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[176].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[176].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[176].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[176].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[176].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[175].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[177].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[177].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[177].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[177].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[177].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[176].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[178].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[178].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[178].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[178].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[178].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[177].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[179].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[179].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[179].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[179].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[179].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[178].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[17].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[17].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[17].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[17].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[17].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[16].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[180].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[180].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[180].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[180].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[180].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[179].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[181].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[181].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[181].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[181].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[181].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[180].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[182].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[182].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[182].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[182].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[182].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[181].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[183].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[183].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[183].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[183].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[183].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[182].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[184].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[184].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[184].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[184].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[184].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[183].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[185].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[185].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[185].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[185].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[185].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[184].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[186].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[186].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[186].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[186].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[186].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[185].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[187].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[187].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[187].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[187].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[187].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[186].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[188].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[188].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[188].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[188].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[188].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[187].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[189].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[189].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[189].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[189].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[189].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[188].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[18].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[18].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[18].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[18].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[18].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[17].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[190].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[190].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[190].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[190].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[190].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[189].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[191].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[191].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[191].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[191].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[191].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[190].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[192].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[192].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[192].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[192].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[192].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[191].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[193].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[193].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[193].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[193].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[193].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[192].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[194].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[194].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[194].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[194].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[194].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[193].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[195].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[195].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[195].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[195].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[195].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[194].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[196].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[196].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[196].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[196].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[196].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[195].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[197].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[197].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[197].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[197].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[197].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[196].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[198].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[198].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[198].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[198].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[198].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[197].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[199].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[199].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[199].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[199].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[199].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[198].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[19].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[19].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[19].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[19].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[19].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[18].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[1].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[1].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[1].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[1].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[1].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[0].genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[200].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[200].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[200].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[200].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[200].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[199].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[201].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[201].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[201].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[201].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[201].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[200].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[202].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[202].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[202].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[202].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[202].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[201].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[203].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[203].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[203].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[203].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[203].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[202].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[204].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[204].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[204].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[204].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[204].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[203].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[205].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[205].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[205].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[205].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[205].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[204].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[206].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[206].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[206].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[206].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[206].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[205].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[207].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[207].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[207].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[207].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[207].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[206].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[208].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[208].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[208].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[208].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[208].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[207].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[209].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[209].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[209].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[209].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[209].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[208].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[20].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[20].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[20].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[20].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[20].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[19].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[210].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[210].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[210].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[210].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[210].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[209].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[211].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[211].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[211].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[211].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[211].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[210].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[212].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[212].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[212].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[212].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[212].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[211].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[213].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[213].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[213].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[213].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[213].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[212].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[214].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[214].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[214].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[214].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[214].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[213].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[215].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[215].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[215].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[215].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[215].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[214].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[216].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[216].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[216].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[216].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[216].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[215].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[217].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[217].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[217].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[217].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[217].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[216].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[218].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[218].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[218].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[218].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[218].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[217].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[219].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[219].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[219].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[219].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[219].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[218].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[21].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[21].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[21].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[21].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[21].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[20].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[220].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[220].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[220].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[220].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[220].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[219].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[221].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[221].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[221].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[221].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[221].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[220].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[222].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[222].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[222].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[222].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[222].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[221].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[223].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[223].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[223].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[223].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[223].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[222].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[224].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[224].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[224].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[224].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[224].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[223].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[225].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[225].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[225].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[225].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[225].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[224].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[226].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[226].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[226].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[226].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[226].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[225].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[227].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[227].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[227].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[227].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[227].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[226].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[228].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[228].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[228].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[228].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[228].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[227].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[229].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[229].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[229].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[229].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[229].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[228].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[22].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[22].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[22].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[22].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[22].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[21].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[230].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[230].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[230].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[230].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[230].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[229].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[231].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[231].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[231].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[231].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[231].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[230].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[232].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[232].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[232].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[232].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[232].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[231].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[233].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[233].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[233].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[233].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[233].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[232].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[234].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[234].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[234].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[234].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[234].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[233].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[235].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[235].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[235].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[235].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[235].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[234].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[236].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[236].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[236].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[236].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[236].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[235].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[237].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[237].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[237].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[237].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[237].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[236].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[238].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[238].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[238].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[238].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[238].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[237].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[239].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[239].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[239].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[239].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[239].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[238].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[23].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[23].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[23].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[23].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[23].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[22].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[240].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[240].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[240].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[240].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[240].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[239].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[241].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[241].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[241].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[241].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[241].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[240].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[242].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[242].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[242].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[242].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[242].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[241].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[243].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[243].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[243].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[243].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[243].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[242].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[244].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[244].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[244].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[244].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[244].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[243].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[245].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[245].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[245].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[245].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[245].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[244].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[246].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[246].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[246].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[246].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[246].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[245].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[247].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[247].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[247].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[247].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[247].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[246].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[248].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[248].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[248].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[248].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[248].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[247].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[249].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[249].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[249].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[249].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[249].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[248].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[24].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[24].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[24].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[24].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[24].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[23].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[250].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[250].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[250].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[250].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[250].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[249].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[251].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[251].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[251].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[251].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[251].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[250].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[252].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[252].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[252].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[252].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[252].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[251].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[253].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[253].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[253].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[253].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[253].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[252].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[254].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[254].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[254].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[254].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[254].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[253].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[255].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[255].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[255].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[255].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[255].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[254].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[256].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[256].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[256].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[256].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[256].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[255].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[257].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[257].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[257].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[257].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[257].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[256].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[258].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[258].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[258].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[258].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[258].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[257].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[259].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[259].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[259].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[259].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[259].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[258].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[25].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[25].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[25].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[25].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[25].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[24].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[260].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[260].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[260].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[260].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[260].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[259].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[261].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[261].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[261].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[261].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[261].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[260].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[262].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[262].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[262].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[262].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[262].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[261].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[263].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[263].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[263].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[263].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[263].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[262].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[264].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[264].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[264].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[264].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[264].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[263].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[265].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[265].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[265].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[265].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[265].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[264].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[266].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[266].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[266].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[266].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[266].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[265].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[267].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[267].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[267].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[267].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[267].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[266].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[268].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[268].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[268].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[268].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[268].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[267].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[269].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[269].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[269].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[269].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[269].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[268].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[26].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[26].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[26].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[26].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[26].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[25].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[270].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[270].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[270].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[270].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[270].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[269].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[271].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[271].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[271].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[271].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[271].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[270].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[272].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[272].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[272].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[272].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[272].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[271].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[273].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[273].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[273].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[273].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[273].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[272].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[274].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[274].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[274].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[274].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[274].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[273].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[275].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[275].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[275].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[275].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[275].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[274].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[276].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[276].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[276].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[276].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[276].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[275].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[277].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[277].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[277].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[277].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[277].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[276].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[278].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[278].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[278].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[278].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[278].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[277].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[279].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[279].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[279].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[279].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[279].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[278].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[27].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[27].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[27].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[27].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[27].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[26].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[280].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[280].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[280].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[280].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[280].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[279].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[281].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[281].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[281].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[281].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[281].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[280].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[282].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[282].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[282].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[282].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[282].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[281].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[283].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[283].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[283].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[283].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[283].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[282].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[284].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[284].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[284].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[284].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[284].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[283].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[285].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[285].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[285].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[285].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[285].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[284].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[286].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[286].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[286].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[286].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[286].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[285].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[287].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[287].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[287].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[287].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[287].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[286].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[288].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[288].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[288].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[288].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[288].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[287].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[289].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[289].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[289].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[289].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[289].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[288].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[28].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[28].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[28].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[28].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[28].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[27].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[290].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[290].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[290].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[290].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[290].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[289].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[291].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[291].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[291].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[291].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[291].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[290].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[292].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[292].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[292].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[292].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[292].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[291].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[293].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[293].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[293].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[293].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[293].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[292].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[294].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[294].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[294].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[294].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[294].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[293].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[295].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[295].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[295].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[295].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[295].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[294].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[296].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[296].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[296].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[296].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[296].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[295].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[297].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[297].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[297].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[297].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[297].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[296].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[298].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[298].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[298].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[298].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[298].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[297].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[299].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[299].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[299].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[299].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[299].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[298].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[29].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[29].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[29].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[29].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[29].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[28].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[2].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[2].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[2].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[2].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[2].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[1].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[300].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[300].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[300].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[300].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[300].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[299].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[301].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[301].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[301].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[301].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[301].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[300].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[302].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[302].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[302].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[302].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[302].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[301].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[303].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[303].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[303].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[303].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[303].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[302].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[304].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[304].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[304].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[304].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[304].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[303].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[305].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[305].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[305].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[305].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[305].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[304].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[306].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[306].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[306].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[306].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[306].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[305].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[307].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[307].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[307].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[307].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[307].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[306].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[308].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[308].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[308].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[308].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[308].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[307].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[309].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[309].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[309].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[309].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[309].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[308].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[30].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[30].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[30].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[30].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[30].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[29].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[310].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[310].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[310].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[310].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[310].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[309].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[311].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[311].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[311].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[311].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[311].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[310].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[312].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[312].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[312].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[312].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[312].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[311].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[313].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[313].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[313].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[313].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[313].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[312].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[314].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[314].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[314].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[314].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[314].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[313].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[315].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[315].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[315].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[315].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[315].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[314].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[316].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[316].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[316].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[316].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[316].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[315].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[317].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[317].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[317].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[317].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[317].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[316].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[318].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[318].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[318].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[318].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[318].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[317].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[319].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[319].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[319].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[319].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[319].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[318].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[31].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[31].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[31].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[31].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[31].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[30].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[320].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[320].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[320].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[320].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[320].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[319].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[321].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[321].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[321].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[321].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[321].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[320].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[322].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[322].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[322].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[322].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[322].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[321].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[323].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[323].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[323].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[323].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[323].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[322].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[324].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[324].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[324].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[324].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[324].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[323].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[325].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[325].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[325].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[325].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[325].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[324].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[326].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[326].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[326].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[326].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[326].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[325].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[327].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[327].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[327].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[327].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[327].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[326].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[328].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[328].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[328].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[328].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[328].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[327].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[329].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[329].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[329].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[329].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[329].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[328].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[32].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[32].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[32].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[32].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[32].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[31].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[330].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[330].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[330].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[330].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[330].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[329].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[331].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[331].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[331].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[331].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[331].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[330].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[332].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[332].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[332].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[332].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[332].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[331].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[333].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[333].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[333].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[333].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[333].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[332].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[334].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[334].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[334].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[334].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[334].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[333].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[335].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[335].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[335].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[335].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[335].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[334].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[336].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[336].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[336].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[336].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[336].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[335].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[337].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[337].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[337].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[337].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[337].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[336].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[338].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[338].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[338].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[338].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[338].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[337].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[339].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[339].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[339].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[339].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[339].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[338].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[33].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[33].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[33].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[33].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[33].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[32].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[340].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[340].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[340].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[340].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[340].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[339].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[341].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[341].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[341].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[341].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[341].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[340].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[342].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[342].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[342].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[342].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[342].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[341].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[343].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[343].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[343].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[343].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[343].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[342].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[344].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[344].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[344].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[344].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[344].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[343].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[345].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[345].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[345].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[345].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[345].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[344].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[346].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[346].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[346].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[346].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[346].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[345].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[347].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[347].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[347].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[347].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[347].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[346].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[348].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[348].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[348].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[348].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[348].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[347].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[349].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[349].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[349].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[349].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[349].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[348].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[34].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[34].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[34].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[34].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[34].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[33].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[350].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[350].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[350].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[350].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[350].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[349].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[351].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[351].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[351].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[351].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[351].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[350].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[352].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[352].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[352].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[352].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[352].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[351].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[353].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[353].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[353].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[353].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[353].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[352].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[354].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[354].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[354].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[354].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[354].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[353].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[355].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[355].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[355].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[355].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[355].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[354].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[356].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[356].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[356].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[356].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[356].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[355].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[357].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[357].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[357].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[357].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[357].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[356].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[358].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[358].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[358].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[358].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[358].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[357].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[359].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[359].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[359].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[359].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[359].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[358].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[35].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[35].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[35].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[35].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[35].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[34].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[360].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[360].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[360].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[360].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[360].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[359].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[361].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[361].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[361].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[361].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[361].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[360].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[362].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[362].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[362].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[362].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[362].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[361].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[363].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[363].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[363].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[363].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[363].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[362].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[364].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[364].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[364].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[364].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[364].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[363].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[365].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[365].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[365].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[365].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[365].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[364].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[366].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[366].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[366].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[366].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[366].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[365].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[367].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[367].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[367].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[367].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[367].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[366].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[368].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[368].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[368].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[368].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[368].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[367].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[369].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[369].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[369].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[369].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[369].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[368].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[36].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[36].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[36].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[36].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[36].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[35].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[370].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[370].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[370].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[370].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[370].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[369].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[371].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[371].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[371].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[371].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[371].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[370].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[372].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[372].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[372].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[372].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[372].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[371].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[373].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[373].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[373].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[373].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[373].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[372].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[374].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[374].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[374].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[374].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[374].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[373].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[375].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[375].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[375].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[375].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[375].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[374].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[376].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[376].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[376].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[376].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[376].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[375].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[377].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[377].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[377].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[377].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[377].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[376].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[378].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[378].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[378].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[378].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[378].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[377].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[379].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[379].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[379].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[379].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[379].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[378].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[37].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[37].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[37].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[37].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[37].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[36].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[380].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[380].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[380].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[380].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[380].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[379].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[381].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[381].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[381].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[381].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[381].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[380].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[382].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[382].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[382].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[382].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[382].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[381].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[383].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[383].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[383].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[383].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[383].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[382].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[384].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[384].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[384].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[384].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[384].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[383].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[385].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[385].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[385].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[385].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[385].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[384].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[386].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[386].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[386].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[386].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[386].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[385].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[387].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[387].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[387].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[387].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[387].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[386].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[388].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[388].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[388].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[388].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[388].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[387].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[389].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[389].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[389].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[389].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[389].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[388].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[38].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[38].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[38].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[38].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[38].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[37].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[390].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[390].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[390].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[390].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[390].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[389].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[391].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[391].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[391].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[391].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[391].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[390].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[392].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[392].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[392].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[392].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[392].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[391].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[393].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[393].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[393].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[393].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[393].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[392].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[394].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[394].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[394].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[394].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[394].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[393].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[395].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[395].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[395].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[395].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[395].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[394].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[396].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[396].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[396].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[396].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[396].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[395].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[397].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[397].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[397].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[397].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[397].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[396].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[398].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[398].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[398].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[398].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[398].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[397].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[399].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[399].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[399].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[399].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[399].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[398].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[39].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[39].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[39].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[39].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[39].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[38].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[3].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[3].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[3].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[3].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[3].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[2].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[400].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[400].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[400].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[400].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[400].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[399].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[401].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[401].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[401].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[401].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[401].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[400].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[402].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[402].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[402].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[402].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[402].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[401].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[403].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[403].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[403].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[403].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[403].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[402].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[404].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[404].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[404].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[404].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[404].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[403].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[405].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[405].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[405].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[405].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[405].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[404].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[406].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[406].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[406].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[406].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[406].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[405].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[407].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[407].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[407].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[407].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[407].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[406].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[408].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[408].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[408].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[408].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[408].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[407].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[409].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[409].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[409].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[409].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[409].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[408].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[40].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[40].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[40].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[40].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[40].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[39].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[410].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[410].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[410].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[410].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[410].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[409].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[411].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[411].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[411].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[411].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[411].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[410].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[412].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[412].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[412].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[412].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[412].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[411].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[413].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[413].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[413].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[413].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[413].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[412].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[414].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[414].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[414].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[414].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[414].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[413].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[415].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[415].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[415].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[415].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[415].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[414].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[416].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[416].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[416].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[416].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[416].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[415].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[417].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[417].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[417].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[417].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[417].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[416].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[418].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[418].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[418].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[418].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[418].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[417].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[419].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[419].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[419].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[419].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[419].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[418].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[41].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[41].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[41].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[41].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[41].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[40].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[420].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[420].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[420].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[420].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[420].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[419].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[421].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[421].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[421].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[421].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[421].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[420].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[422].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[422].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[422].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[422].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[422].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[421].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[423].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[423].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[423].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[423].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[423].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[422].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[424].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[424].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[424].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[424].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[424].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[423].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[425].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[425].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[425].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[425].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[425].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[424].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[426].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[426].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[426].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[426].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[426].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[425].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[427].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[427].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[427].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[427].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[427].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[426].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[428].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[428].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[428].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[428].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[428].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[427].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[429].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[429].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[429].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[429].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[429].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[428].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[42].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[42].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[42].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[42].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[42].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[41].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[430].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[430].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[430].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[430].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[430].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[429].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[431].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[431].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[431].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[431].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[431].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[430].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[432].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[432].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[432].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[432].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[432].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[431].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[433].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[433].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[433].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[433].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[433].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[432].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[434].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[434].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[434].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[434].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[434].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[433].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[435].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[435].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[435].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[435].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[435].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[434].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[436].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[436].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[436].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[436].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[436].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[435].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[437].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[437].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[437].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[437].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[437].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[436].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[438].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[438].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[438].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[438].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[438].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[437].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[439].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[439].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[439].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[439].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[439].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[438].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[43].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[43].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[43].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[43].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[43].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[42].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[440].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[440].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[440].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[440].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[440].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[439].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[441].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[441].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[441].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[441].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[441].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[440].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[442].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[442].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[442].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[442].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[442].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[441].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[443].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[443].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[443].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[443].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[443].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[442].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[444].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[444].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[444].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[444].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[444].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[443].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[445].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[445].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[445].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[445].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[445].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[444].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[446].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[446].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[446].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[446].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[446].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[445].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[447].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[447].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[447].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[447].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[447].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[446].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[448].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[448].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[448].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[448].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[448].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[447].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[449].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[449].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[449].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[449].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[449].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[448].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[44].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[44].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[44].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[44].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[44].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[43].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[450].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[450].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[450].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[450].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[450].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[449].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[451].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[451].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[451].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[451].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[451].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[450].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[452].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[452].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[452].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[452].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[452].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[451].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[453].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[453].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[453].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[453].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[453].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[452].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[454].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[454].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[454].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[454].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[454].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[453].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[455].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[455].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[455].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[455].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[455].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[454].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[456].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[456].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[456].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[456].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[456].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[455].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[457].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[457].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[457].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[457].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[457].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[456].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[458].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[458].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[458].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[458].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[458].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[457].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[459].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[459].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[459].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[459].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[459].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[458].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[45].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[45].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[45].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[45].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[45].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[44].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[460].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[460].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[460].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[460].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[460].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[459].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[461].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[461].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[461].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[461].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[461].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[460].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[462].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[462].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[462].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[462].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[462].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[461].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[463].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[463].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[463].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[463].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[463].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[462].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[464].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[464].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[464].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[464].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[464].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[463].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[465].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[465].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[465].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[465].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[465].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[464].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[466].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[466].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[466].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[466].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[466].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[465].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[467].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[467].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[467].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[467].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[467].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[466].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[468].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[468].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[468].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[468].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[468].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[467].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[469].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[469].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[469].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[469].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[469].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[468].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[46].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[46].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[46].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[46].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[46].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[45].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[470].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[470].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[470].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[470].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[470].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[469].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[471].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[471].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[471].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[471].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[471].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[470].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[472].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[472].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[472].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[472].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[472].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[471].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[473].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[473].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[473].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[473].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[473].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[472].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[474].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[474].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[474].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[474].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[474].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[473].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[475].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[475].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[475].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[475].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[475].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[474].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[476].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[476].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[476].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[476].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[476].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[475].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[477].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[477].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[477].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[477].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[477].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[476].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[478].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[478].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[478].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[478].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[478].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[477].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[479].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[479].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[479].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[479].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[479].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[478].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[47].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[47].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[47].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[47].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[47].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[46].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[480].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[480].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[480].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[480].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[480].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[479].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[481].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[481].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[481].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[481].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[481].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[480].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[482].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[482].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[482].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[482].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[482].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[481].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[483].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[483].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[483].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[483].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[483].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[482].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[484].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[484].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[484].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[484].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[484].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[483].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[485].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[485].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[485].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[485].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[485].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[484].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[486].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[486].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[486].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[486].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[486].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[485].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[487].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[487].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[487].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[487].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[487].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[486].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[488].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[488].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[488].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[488].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[488].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[487].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[489].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[489].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[489].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[489].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[489].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[488].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[48].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[48].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[48].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[48].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[48].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[47].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[490].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[490].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[490].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[490].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[490].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[489].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[491].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[491].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[491].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[491].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[491].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[490].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[492].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[492].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[492].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[492].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[492].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[491].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[493].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[493].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[493].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[493].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[493].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[492].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[494].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[494].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[494].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[494].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[494].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[493].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[495].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[495].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[495].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[495].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[495].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[494].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[496].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[496].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[496].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[496].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[496].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[495].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[497].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[497].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[497].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[497].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[497].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[496].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[498].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[498].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[498].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[498].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[498].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[497].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[499].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[499].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[499].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[499].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[499].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[498].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[49].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[49].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[49].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[49].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[49].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[48].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[4].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[4].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[4].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[4].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[4].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[3].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[500].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[500].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[500].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[500].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[500].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[499].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[501].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[501].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[501].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[501].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[501].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[500].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[502].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[502].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[502].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[502].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[502].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[501].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[503].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[503].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[503].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[503].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[503].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[502].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[504].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[504].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[504].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[504].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[504].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[503].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[505].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[505].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[505].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[505].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[505].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[504].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[506].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[506].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[506].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[506].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[506].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[505].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[507].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[507].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[507].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[507].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[507].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[506].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[508].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[508].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[508].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[508].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[508].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[507].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[509].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[509].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[509].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[509].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[509].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[508].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[50].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[50].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[50].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[50].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[50].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[49].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[510].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[510].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[510].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[510].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[510].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[509].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[511].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[511].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[511].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[511].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[511].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[510].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[51].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[51].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[51].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[51].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[51].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[50].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[52].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[52].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[52].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[52].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[52].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[51].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[53].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[53].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[53].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[53].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[53].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[52].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[54].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[54].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[54].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[54].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[54].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[53].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[55].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[55].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[55].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[55].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[55].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[54].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[56].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[56].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[56].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[56].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[56].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[55].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[57].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[57].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[57].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[57].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[57].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[56].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[58].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[58].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[58].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[58].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[58].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[57].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[59].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[59].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[59].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[59].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[59].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[58].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[5].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[5].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[5].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[5].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[5].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[4].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[60].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[60].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[60].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[60].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[60].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[59].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[61].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[61].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[61].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[61].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[61].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[60].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[62].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[62].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[62].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[62].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[62].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[61].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[63].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[63].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[63].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[63].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[63].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[62].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[64].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[64].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[64].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[64].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[64].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[63].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[65].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[65].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[65].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[65].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[65].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[64].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[66].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[66].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[66].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[66].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[66].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[65].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[67].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[67].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[67].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[67].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[67].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[66].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[68].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[68].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[68].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[68].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[68].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[67].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[69].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[69].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[69].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[69].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[69].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[68].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[6].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[6].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[6].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[6].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[6].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[5].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[70].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[70].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[70].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[70].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[70].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[69].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[71].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[71].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[71].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[71].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[71].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[70].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[72].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[72].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[72].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[72].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[72].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[71].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[73].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[73].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[73].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[73].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[73].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[72].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[74].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[74].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[74].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[74].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[74].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[73].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[75].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[75].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[75].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[75].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[75].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[74].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[76].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[76].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[76].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[76].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[76].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[75].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[77].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[77].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[77].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[77].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[77].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[76].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[78].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[78].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[78].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[78].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[78].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[77].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[79].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[79].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[79].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[79].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[79].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[78].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[7].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[7].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[7].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[7].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[7].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[6].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[80].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[80].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[80].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[80].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[80].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[79].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[81].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[81].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[81].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[81].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[81].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[80].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[82].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[82].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[82].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[82].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[82].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[81].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[83].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[83].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[83].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[83].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[83].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[82].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[84].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[84].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[84].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[84].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[84].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[83].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[85].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[85].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[85].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[85].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[85].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[84].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[86].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[86].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[86].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[86].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[86].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[85].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[87].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[87].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[87].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[87].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[87].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[86].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[88].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[88].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[88].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[88].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[88].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[87].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[89].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[89].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[89].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[89].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[89].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[88].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[8].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[8].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[8].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[8].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[8].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[7].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[90].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[90].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[90].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[90].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[90].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[89].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[91].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[91].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[91].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[91].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[91].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[90].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[92].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[92].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[92].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[92].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[92].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[91].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[93].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[93].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[93].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[93].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[93].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[92].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[94].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[94].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[94].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[94].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[94].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[93].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[95].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[95].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[95].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[95].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[95].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[94].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[96].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[96].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[96].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[96].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[96].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[95].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[97].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[97].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[97].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[97].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[97].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[96].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[98].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[98].genblk1.genblk1.latch.clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[98].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[98].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[98].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[97].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[99].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[100].genblk1.genblk1.latch.clkout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[99].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[99].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[99].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[98].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[9].genblk1.genblk1.latch.u_inv1.inv  (.A(\shift_reg[10].genblk1.genblk1.latch.clkout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[9].genblk1.genblk1.latch.nclk ));
 sky130_fd_sc_hd__inv_1 \shift_reg[9].genblk1.genblk1.latch.u_inv2.inv  (.A(\shift_reg[9].genblk1.genblk1.latch.nclk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\shift_reg[8].genblk1.genblk1.latch.clk ));
 sky130_fd_sc_hd__inv_1 \u_invA.inv  (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_invA.out ));
 sky130_fd_sc_hd__inv_1 \u_invB.inv  (.A(\u_invA.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_invB.out ));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__conb_1 _513__3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net3));
 sky130_fd_sc_hd__conb_1 _514__4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net4));
 sky130_fd_sc_hd__conb_1 _515__5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net5));
 sky130_fd_sc_hd__conb_1 _516__6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net6));
 sky130_fd_sc_hd__conb_1 _517__7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net7));
 sky130_fd_sc_hd__conb_1 _518__8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net8));
 sky130_fd_sc_hd__conb_1 _519__9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net9));
 sky130_fd_sc_hd__conb_1 _520__10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__conb_1 _521__11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net11));
 sky130_fd_sc_hd__conb_1 _522__12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net12));
 sky130_fd_sc_hd__conb_1 _523__13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net13));
 sky130_fd_sc_hd__conb_1 _524__14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net14));
 sky130_fd_sc_hd__conb_1 _525__15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net15));
 sky130_fd_sc_hd__conb_1 _526__16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net16));
 sky130_fd_sc_hd__conb_1 _527__17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net17));
 sky130_fd_sc_hd__conb_1 _528__18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net18));
 sky130_fd_sc_hd__conb_1 _530__19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net19));
 sky130_fd_sc_hd__conb_1 _531__20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__conb_1 _532__21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__conb_1 _533__22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__conb_1 _534__23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net23));
 sky130_fd_sc_hd__conb_1 _535__24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net24));
 sky130_fd_sc_hd__conb_1 _536__25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net25));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_257 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_311 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_86 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_229 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_166 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_308 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
