VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rburt16_bias_generator
  CLASS BLOCK ;
  FOREIGN tt_um_rburt16_bias_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 18.559999 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 780.947205 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 16.850 207.240 19.810 207.245 ;
        RECT 6.020 197.400 11.410 207.240 ;
      LAYER pwell ;
        RECT 11.420 197.400 14.380 207.190 ;
      LAYER nwell ;
        RECT 14.420 197.405 19.810 207.240 ;
      LAYER pwell ;
        RECT 19.830 197.415 22.790 207.205 ;
      LAYER nwell ;
        RECT 22.820 202.660 32.975 207.240 ;
        RECT 35.000 206.000 40.840 208.460 ;
      LAYER pwell ;
        RECT 33.020 202.700 42.980 204.910 ;
      LAYER nwell ;
        RECT 22.820 200.400 42.480 202.660 ;
        RECT 14.420 197.400 17.380 197.405 ;
        RECT 22.820 197.400 32.975 200.400 ;
      LAYER pwell ;
        RECT 33.020 197.400 42.810 200.360 ;
        RECT 6.000 196.990 28.400 197.090 ;
        RECT 6.000 194.200 42.980 196.990 ;
        RECT 6.000 187.300 37.880 194.200 ;
      LAYER nwell ;
        RECT 16.850 181.240 19.810 181.245 ;
        RECT 6.020 171.400 11.410 181.240 ;
      LAYER pwell ;
        RECT 11.420 171.400 14.380 181.190 ;
      LAYER nwell ;
        RECT 14.420 171.405 19.810 181.240 ;
      LAYER pwell ;
        RECT 19.830 171.415 22.790 181.205 ;
      LAYER nwell ;
        RECT 22.820 176.660 32.975 181.240 ;
        RECT 35.000 180.000 40.840 182.460 ;
      LAYER pwell ;
        RECT 33.020 176.700 42.980 178.910 ;
      LAYER nwell ;
        RECT 22.820 174.400 42.480 176.660 ;
        RECT 14.420 171.400 17.380 171.405 ;
        RECT 22.820 171.400 32.975 174.400 ;
      LAYER pwell ;
        RECT 33.020 171.400 42.810 174.360 ;
        RECT 6.000 170.990 28.400 171.090 ;
        RECT 6.000 168.200 42.980 170.990 ;
        RECT 6.000 161.300 37.880 168.200 ;
      LAYER nwell ;
        RECT 16.850 155.240 19.810 155.245 ;
        RECT 6.020 145.400 11.410 155.240 ;
      LAYER pwell ;
        RECT 11.420 145.400 14.380 155.190 ;
      LAYER nwell ;
        RECT 14.420 145.405 19.810 155.240 ;
      LAYER pwell ;
        RECT 19.830 145.415 22.790 155.205 ;
      LAYER nwell ;
        RECT 22.820 150.660 32.975 155.240 ;
        RECT 35.000 154.000 40.840 156.460 ;
      LAYER pwell ;
        RECT 33.020 150.700 42.980 152.910 ;
      LAYER nwell ;
        RECT 22.820 148.400 42.480 150.660 ;
        RECT 14.420 145.400 17.380 145.405 ;
        RECT 22.820 145.400 32.975 148.400 ;
      LAYER pwell ;
        RECT 33.020 145.400 42.810 148.360 ;
        RECT 48.300 146.320 58.090 168.720 ;
      LAYER nwell ;
        RECT 58.400 163.310 68.240 168.700 ;
      LAYER pwell ;
        RECT 58.400 160.340 68.190 163.300 ;
      LAYER nwell ;
        RECT 58.400 157.870 68.240 160.300 ;
        RECT 58.400 157.340 68.245 157.870 ;
        RECT 58.405 154.910 68.245 157.340 ;
      LAYER pwell ;
        RECT 58.415 151.930 68.205 154.890 ;
        RECT 6.000 144.990 28.400 145.090 ;
        RECT 6.000 142.200 42.980 144.990 ;
        RECT 6.000 135.300 37.880 142.200 ;
        RECT 48.300 136.840 57.990 146.320 ;
      LAYER nwell ;
        RECT 58.400 141.745 68.240 151.900 ;
      LAYER pwell ;
        RECT 74.300 146.320 84.090 168.720 ;
      LAYER nwell ;
        RECT 84.400 163.310 94.240 168.700 ;
      LAYER pwell ;
        RECT 84.400 160.340 94.190 163.300 ;
      LAYER nwell ;
        RECT 84.400 157.870 94.240 160.300 ;
        RECT 84.400 157.340 94.245 157.870 ;
        RECT 84.405 154.910 94.245 157.340 ;
      LAYER pwell ;
        RECT 84.415 151.930 94.205 154.890 ;
        RECT 55.200 131.740 57.990 136.840 ;
        RECT 58.400 131.910 61.360 141.700 ;
      LAYER nwell ;
        RECT 61.400 132.240 63.660 141.745 ;
      LAYER pwell ;
        RECT 63.700 131.740 65.910 141.700 ;
      LAYER nwell ;
        RECT 67.000 134.000 69.460 139.840 ;
      LAYER pwell ;
        RECT 74.300 136.840 83.990 146.320 ;
      LAYER nwell ;
        RECT 84.400 141.745 94.240 151.900 ;
      LAYER pwell ;
        RECT 81.200 131.740 83.990 136.840 ;
        RECT 84.400 131.910 87.360 141.700 ;
      LAYER nwell ;
        RECT 87.400 132.240 89.660 141.745 ;
      LAYER pwell ;
        RECT 89.700 131.740 91.910 141.700 ;
      LAYER nwell ;
        RECT 93.000 134.000 95.460 139.840 ;
        RECT 16.850 129.240 19.810 129.245 ;
        RECT 6.020 119.400 11.410 129.240 ;
      LAYER pwell ;
        RECT 11.420 119.400 14.380 129.190 ;
      LAYER nwell ;
        RECT 14.420 119.405 19.810 129.240 ;
      LAYER pwell ;
        RECT 19.830 119.415 22.790 129.205 ;
      LAYER nwell ;
        RECT 22.820 124.660 32.975 129.240 ;
        RECT 35.000 128.000 40.840 130.460 ;
      LAYER pwell ;
        RECT 33.020 124.700 42.980 126.910 ;
      LAYER nwell ;
        RECT 22.820 122.400 42.480 124.660 ;
        RECT 14.420 119.400 17.380 119.405 ;
        RECT 22.820 119.400 32.975 122.400 ;
      LAYER pwell ;
        RECT 33.020 119.400 42.810 122.360 ;
        RECT 6.000 118.990 28.400 119.090 ;
        RECT 6.000 116.200 42.980 118.990 ;
        RECT 6.000 109.300 37.880 116.200 ;
      LAYER nwell ;
        RECT 16.850 103.240 19.810 103.245 ;
        RECT 6.020 93.400 11.410 103.240 ;
      LAYER pwell ;
        RECT 11.420 93.400 14.380 103.190 ;
      LAYER nwell ;
        RECT 14.420 93.405 19.810 103.240 ;
      LAYER pwell ;
        RECT 19.830 93.415 22.790 103.205 ;
      LAYER nwell ;
        RECT 22.820 98.660 32.975 103.240 ;
        RECT 35.000 102.000 40.840 104.460 ;
      LAYER pwell ;
        RECT 48.300 104.320 58.090 126.720 ;
      LAYER nwell ;
        RECT 58.400 121.310 68.240 126.700 ;
      LAYER pwell ;
        RECT 58.400 118.340 68.190 121.300 ;
      LAYER nwell ;
        RECT 58.400 115.870 68.240 118.300 ;
        RECT 58.400 115.340 68.245 115.870 ;
        RECT 58.405 112.910 68.245 115.340 ;
      LAYER pwell ;
        RECT 58.415 109.930 68.205 112.890 ;
        RECT 33.020 98.700 42.980 100.910 ;
      LAYER nwell ;
        RECT 22.820 96.400 42.480 98.660 ;
        RECT 14.420 93.400 17.380 93.405 ;
        RECT 22.820 93.400 32.975 96.400 ;
      LAYER pwell ;
        RECT 33.020 93.400 42.810 96.360 ;
        RECT 48.300 94.840 57.990 104.320 ;
      LAYER nwell ;
        RECT 58.400 99.745 68.240 109.900 ;
      LAYER pwell ;
        RECT 74.300 104.320 84.090 126.720 ;
      LAYER nwell ;
        RECT 84.400 121.310 94.240 126.700 ;
      LAYER pwell ;
        RECT 84.400 118.340 94.190 121.300 ;
      LAYER nwell ;
        RECT 84.400 115.870 94.240 118.300 ;
        RECT 84.400 115.340 94.245 115.870 ;
        RECT 84.405 112.910 94.245 115.340 ;
      LAYER pwell ;
        RECT 84.415 109.930 94.205 112.890 ;
        RECT 6.000 92.990 28.400 93.090 ;
        RECT 6.000 90.200 42.980 92.990 ;
        RECT 6.000 83.300 37.880 90.200 ;
        RECT 55.200 89.740 57.990 94.840 ;
        RECT 58.400 89.910 61.360 99.700 ;
      LAYER nwell ;
        RECT 61.400 90.240 63.660 99.745 ;
      LAYER pwell ;
        RECT 63.700 89.740 65.910 99.700 ;
      LAYER nwell ;
        RECT 67.000 92.000 69.460 97.840 ;
      LAYER pwell ;
        RECT 74.300 94.840 83.990 104.320 ;
      LAYER nwell ;
        RECT 84.400 99.745 94.240 109.900 ;
      LAYER pwell ;
        RECT 81.200 89.740 83.990 94.840 ;
        RECT 84.400 89.910 87.360 99.700 ;
      LAYER nwell ;
        RECT 87.400 90.240 89.660 99.745 ;
      LAYER pwell ;
        RECT 89.700 89.740 91.910 99.700 ;
      LAYER nwell ;
        RECT 93.000 92.000 95.460 97.840 ;
        RECT 16.850 77.240 19.810 77.245 ;
        RECT 6.020 67.400 11.410 77.240 ;
      LAYER pwell ;
        RECT 11.420 67.400 14.380 77.190 ;
      LAYER nwell ;
        RECT 14.420 67.405 19.810 77.240 ;
      LAYER pwell ;
        RECT 19.830 67.415 22.790 77.205 ;
      LAYER nwell ;
        RECT 22.820 72.660 32.975 77.240 ;
        RECT 35.000 76.000 40.840 78.460 ;
      LAYER pwell ;
        RECT 33.020 72.700 42.980 74.910 ;
      LAYER nwell ;
        RECT 22.820 70.400 42.480 72.660 ;
        RECT 14.420 67.400 17.380 67.405 ;
        RECT 22.820 67.400 32.975 70.400 ;
      LAYER pwell ;
        RECT 33.020 67.400 42.810 70.360 ;
        RECT 6.000 66.990 28.400 67.090 ;
        RECT 6.000 64.200 42.980 66.990 ;
        RECT 6.000 57.300 37.880 64.200 ;
        RECT 48.300 62.320 58.090 84.720 ;
      LAYER nwell ;
        RECT 58.400 79.310 68.240 84.700 ;
      LAYER pwell ;
        RECT 58.400 76.340 68.190 79.300 ;
      LAYER nwell ;
        RECT 58.400 73.870 68.240 76.300 ;
        RECT 58.400 73.340 68.245 73.870 ;
        RECT 58.405 70.910 68.245 73.340 ;
      LAYER pwell ;
        RECT 58.415 67.930 68.205 70.890 ;
        RECT 48.300 52.840 57.990 62.320 ;
      LAYER nwell ;
        RECT 58.400 57.745 68.240 67.900 ;
      LAYER pwell ;
        RECT 74.300 62.320 84.090 84.720 ;
      LAYER nwell ;
        RECT 84.400 79.310 94.240 84.700 ;
      LAYER pwell ;
        RECT 84.400 76.340 94.190 79.300 ;
      LAYER nwell ;
        RECT 84.400 73.870 94.240 76.300 ;
        RECT 84.400 73.340 94.245 73.870 ;
        RECT 84.405 70.910 94.245 73.340 ;
      LAYER pwell ;
        RECT 84.415 67.930 94.205 70.890 ;
      LAYER nwell ;
        RECT 16.850 51.240 19.810 51.245 ;
        RECT 6.020 41.400 11.410 51.240 ;
      LAYER pwell ;
        RECT 11.420 41.400 14.380 51.190 ;
      LAYER nwell ;
        RECT 14.420 41.405 19.810 51.240 ;
      LAYER pwell ;
        RECT 19.830 41.415 22.790 51.205 ;
      LAYER nwell ;
        RECT 22.820 46.660 32.975 51.240 ;
        RECT 35.000 50.000 40.840 52.460 ;
      LAYER pwell ;
        RECT 33.020 46.700 42.980 48.910 ;
        RECT 55.200 47.740 57.990 52.840 ;
        RECT 58.400 47.910 61.360 57.700 ;
      LAYER nwell ;
        RECT 61.400 48.240 63.660 57.745 ;
      LAYER pwell ;
        RECT 63.700 47.740 65.910 57.700 ;
      LAYER nwell ;
        RECT 67.000 50.000 69.460 55.840 ;
      LAYER pwell ;
        RECT 74.300 52.840 83.990 62.320 ;
      LAYER nwell ;
        RECT 84.400 57.745 94.240 67.900 ;
      LAYER pwell ;
        RECT 81.200 47.740 83.990 52.840 ;
        RECT 84.400 47.910 87.360 57.700 ;
      LAYER nwell ;
        RECT 87.400 48.240 89.660 57.745 ;
      LAYER pwell ;
        RECT 89.700 47.740 91.910 57.700 ;
      LAYER nwell ;
        RECT 93.000 50.000 95.460 55.840 ;
        RECT 22.820 44.400 42.480 46.660 ;
        RECT 14.420 41.400 17.380 41.405 ;
        RECT 22.820 41.400 32.975 44.400 ;
      LAYER pwell ;
        RECT 33.020 41.400 42.810 44.360 ;
        RECT 6.000 40.990 28.400 41.090 ;
        RECT 6.000 38.200 42.980 40.990 ;
        RECT 6.000 31.300 37.880 38.200 ;
      LAYER nwell ;
        RECT 16.850 25.240 19.810 25.245 ;
        RECT 6.020 15.400 11.410 25.240 ;
      LAYER pwell ;
        RECT 11.420 15.400 14.380 25.190 ;
      LAYER nwell ;
        RECT 14.420 15.405 19.810 25.240 ;
      LAYER pwell ;
        RECT 19.830 15.415 22.790 25.205 ;
      LAYER nwell ;
        RECT 22.820 20.660 32.975 25.240 ;
        RECT 35.000 24.000 40.840 26.460 ;
      LAYER pwell ;
        RECT 33.020 20.700 42.980 22.910 ;
      LAYER nwell ;
        RECT 22.820 18.400 42.480 20.660 ;
      LAYER pwell ;
        RECT 48.300 20.320 58.090 42.720 ;
      LAYER nwell ;
        RECT 58.400 37.310 68.240 42.700 ;
      LAYER pwell ;
        RECT 58.400 34.340 68.190 37.300 ;
      LAYER nwell ;
        RECT 58.400 31.870 68.240 34.300 ;
        RECT 58.400 31.340 68.245 31.870 ;
        RECT 58.405 28.910 68.245 31.340 ;
      LAYER pwell ;
        RECT 58.415 25.930 68.205 28.890 ;
      LAYER nwell ;
        RECT 14.420 15.400 17.380 15.405 ;
        RECT 22.820 15.400 32.975 18.400 ;
      LAYER pwell ;
        RECT 33.020 15.400 42.810 18.360 ;
        RECT 6.000 14.990 28.400 15.090 ;
        RECT 6.000 12.200 42.980 14.990 ;
        RECT 6.000 5.300 37.880 12.200 ;
        RECT 48.300 10.840 57.990 20.320 ;
      LAYER nwell ;
        RECT 58.400 15.745 68.240 25.900 ;
      LAYER pwell ;
        RECT 74.300 20.320 84.090 42.720 ;
      LAYER nwell ;
        RECT 84.400 37.310 94.240 42.700 ;
      LAYER pwell ;
        RECT 84.400 34.340 94.190 37.300 ;
      LAYER nwell ;
        RECT 84.400 31.870 94.240 34.300 ;
        RECT 84.400 31.340 94.245 31.870 ;
        RECT 84.405 28.910 94.245 31.340 ;
      LAYER pwell ;
        RECT 84.415 25.930 94.205 28.890 ;
        RECT 55.200 5.740 57.990 10.840 ;
        RECT 58.400 5.910 61.360 15.700 ;
      LAYER nwell ;
        RECT 61.400 6.240 63.660 15.745 ;
      LAYER pwell ;
        RECT 63.700 5.740 65.910 15.700 ;
      LAYER nwell ;
        RECT 67.000 8.000 69.460 13.840 ;
      LAYER pwell ;
        RECT 74.300 10.840 83.990 20.320 ;
      LAYER nwell ;
        RECT 84.400 15.745 94.240 25.900 ;
      LAYER pwell ;
        RECT 81.200 5.740 83.990 10.840 ;
        RECT 84.400 5.910 87.360 15.700 ;
      LAYER nwell ;
        RECT 87.400 6.240 89.660 15.745 ;
      LAYER pwell ;
        RECT 89.700 5.740 91.910 15.700 ;
      LAYER nwell ;
        RECT 93.000 8.000 95.460 13.840 ;
      LAYER li1 ;
        RECT 35.180 208.110 40.660 208.280 ;
        RECT 17.030 207.060 19.630 207.065 ;
        RECT 6.200 206.890 11.230 207.060 ;
        RECT 6.200 197.750 6.370 206.890 ;
        RECT 7.000 206.375 8.000 206.545 ;
        RECT 6.770 198.120 6.940 206.160 ;
        RECT 8.060 198.120 8.230 206.160 ;
        RECT 8.630 197.750 8.800 206.890 ;
        RECT 9.430 206.375 10.430 206.545 ;
        RECT 9.200 198.120 9.370 206.160 ;
        RECT 10.490 198.120 10.660 206.160 ;
        RECT 11.060 197.750 11.230 206.890 ;
        RECT 6.200 197.580 11.230 197.750 ;
        RECT 11.600 206.840 14.200 207.010 ;
        RECT 11.600 197.750 11.770 206.840 ;
        RECT 12.400 206.330 13.400 206.500 ;
        RECT 12.170 198.120 12.340 206.160 ;
        RECT 13.460 198.120 13.630 206.160 ;
        RECT 14.030 197.750 14.200 206.840 ;
        RECT 11.600 197.580 14.200 197.750 ;
        RECT 14.600 206.895 19.630 207.060 ;
        RECT 14.600 206.890 17.200 206.895 ;
        RECT 14.600 197.750 14.770 206.890 ;
        RECT 15.400 206.375 16.400 206.545 ;
        RECT 15.170 198.120 15.340 206.160 ;
        RECT 16.460 198.120 16.630 206.160 ;
        RECT 17.030 197.755 17.200 206.890 ;
        RECT 17.830 206.380 18.830 206.550 ;
        RECT 17.600 198.125 17.770 206.165 ;
        RECT 18.890 198.125 19.060 206.165 ;
        RECT 19.460 197.755 19.630 206.895 ;
        RECT 17.030 197.750 19.630 197.755 ;
        RECT 14.600 197.585 19.630 197.750 ;
        RECT 20.010 206.855 22.610 207.025 ;
        RECT 20.010 197.765 20.180 206.855 ;
        RECT 20.810 206.345 21.810 206.515 ;
        RECT 20.580 198.135 20.750 206.175 ;
        RECT 21.870 198.135 22.040 206.175 ;
        RECT 22.440 197.765 22.610 206.855 ;
        RECT 20.010 197.595 22.610 197.765 ;
        RECT 23.000 206.890 32.795 207.060 ;
        RECT 23.000 197.750 23.170 206.890 ;
        RECT 23.800 206.375 24.800 206.545 ;
        RECT 23.570 198.120 23.740 206.160 ;
        RECT 24.860 198.120 25.030 206.160 ;
        RECT 25.400 197.750 25.600 206.890 ;
        RECT 26.200 206.375 27.200 206.545 ;
        RECT 25.970 198.120 26.140 206.160 ;
        RECT 27.260 198.120 27.430 206.160 ;
        RECT 27.800 197.750 28.000 206.890 ;
        RECT 28.600 206.375 29.600 206.545 ;
        RECT 28.370 198.120 28.540 206.160 ;
        RECT 29.660 198.120 29.830 206.160 ;
        RECT 30.195 197.750 30.400 206.890 ;
        RECT 30.995 206.375 31.995 206.545 ;
        RECT 30.765 198.120 30.935 206.160 ;
        RECT 32.055 198.120 32.225 206.160 ;
        RECT 32.625 202.480 32.795 206.890 ;
        RECT 35.180 206.350 35.350 208.110 ;
        RECT 35.720 207.540 39.760 207.710 ;
        RECT 39.975 206.980 40.145 207.480 ;
        RECT 35.720 206.750 39.760 206.920 ;
        RECT 40.490 206.350 40.660 208.110 ;
        RECT 35.180 206.180 40.660 206.350 ;
        RECT 33.200 204.560 42.800 204.730 ;
        RECT 33.200 203.050 33.370 204.560 ;
        RECT 34.000 204.050 42.000 204.220 ;
        RECT 33.770 203.420 33.940 203.880 ;
        RECT 42.060 203.420 42.230 203.880 ;
        RECT 42.630 203.050 42.800 204.560 ;
        RECT 33.200 202.880 42.800 203.050 ;
        RECT 32.625 202.310 42.300 202.480 ;
        RECT 32.625 200.750 32.870 202.310 ;
        RECT 33.500 201.795 41.500 201.965 ;
        RECT 33.270 201.120 33.440 201.580 ;
        RECT 41.560 201.120 41.730 201.580 ;
        RECT 42.130 200.750 42.300 202.310 ;
        RECT 32.625 200.580 42.300 200.750 ;
        RECT 32.625 197.750 32.795 200.580 ;
        RECT 14.600 197.580 17.200 197.585 ;
        RECT 23.000 197.580 32.795 197.750 ;
        RECT 33.200 200.010 42.630 200.180 ;
        RECT 33.200 197.750 33.370 200.010 ;
        RECT 33.740 199.440 41.780 199.610 ;
        RECT 41.950 198.380 42.120 199.380 ;
        RECT 33.740 198.150 41.780 198.320 ;
        RECT 42.460 197.750 42.630 200.010 ;
        RECT 33.200 197.580 42.630 197.750 ;
        RECT 6.180 196.810 28.220 196.910 ;
        RECT 6.180 196.740 42.800 196.810 ;
        RECT 6.180 187.650 6.350 196.740 ;
        RECT 6.980 196.230 7.980 196.400 ;
        RECT 6.750 188.020 6.920 196.060 ;
        RECT 8.040 188.020 8.210 196.060 ;
        RECT 8.610 187.650 8.780 196.740 ;
        RECT 9.410 196.230 10.410 196.400 ;
        RECT 9.180 188.020 9.350 196.060 ;
        RECT 10.470 188.020 10.640 196.060 ;
        RECT 11.040 187.650 11.210 196.740 ;
        RECT 11.840 196.230 12.840 196.400 ;
        RECT 11.610 188.020 11.780 196.060 ;
        RECT 12.900 188.020 13.070 196.060 ;
        RECT 13.470 187.650 13.640 196.740 ;
        RECT 14.270 196.230 15.270 196.400 ;
        RECT 14.040 188.020 14.210 196.060 ;
        RECT 15.330 188.020 15.500 196.060 ;
        RECT 15.900 187.650 16.070 196.740 ;
        RECT 16.700 196.230 17.700 196.400 ;
        RECT 16.470 188.020 16.640 196.060 ;
        RECT 17.760 188.020 17.930 196.060 ;
        RECT 18.330 187.650 18.500 196.740 ;
        RECT 19.130 196.230 20.130 196.400 ;
        RECT 18.900 188.020 19.070 196.060 ;
        RECT 20.190 188.020 20.360 196.060 ;
        RECT 20.760 187.650 20.930 196.740 ;
        RECT 21.560 196.230 22.560 196.400 ;
        RECT 21.330 188.020 21.500 196.060 ;
        RECT 22.620 188.020 22.790 196.060 ;
        RECT 23.190 187.650 23.360 196.740 ;
        RECT 23.990 196.230 24.990 196.400 ;
        RECT 23.760 188.020 23.930 196.060 ;
        RECT 25.050 188.020 25.220 196.060 ;
        RECT 25.620 187.650 25.790 196.740 ;
        RECT 28.050 196.640 42.800 196.740 ;
        RECT 26.420 196.230 27.420 196.400 ;
        RECT 26.190 188.020 26.360 196.060 ;
        RECT 27.480 188.020 27.650 196.060 ;
        RECT 28.050 194.550 28.270 196.640 ;
        RECT 28.900 196.130 42.000 196.300 ;
        RECT 28.670 194.920 28.840 195.960 ;
        RECT 42.060 194.920 42.230 195.960 ;
        RECT 42.630 194.550 42.800 196.640 ;
        RECT 28.050 194.380 42.800 194.550 ;
        RECT 28.050 194.340 37.700 194.380 ;
        RECT 28.050 192.250 28.270 194.340 ;
        RECT 28.900 193.830 36.900 194.000 ;
        RECT 28.670 192.620 28.840 193.660 ;
        RECT 36.960 192.620 37.130 193.660 ;
        RECT 37.530 192.250 37.700 194.340 ;
        RECT 28.050 192.040 37.700 192.250 ;
        RECT 28.050 189.950 28.270 192.040 ;
        RECT 28.900 191.530 36.900 191.700 ;
        RECT 28.670 190.320 28.840 191.360 ;
        RECT 36.960 190.320 37.130 191.360 ;
        RECT 37.530 189.950 37.700 192.040 ;
        RECT 28.050 189.740 37.700 189.950 ;
        RECT 28.050 187.650 28.270 189.740 ;
        RECT 28.900 189.230 36.900 189.400 ;
        RECT 28.670 188.020 28.840 189.060 ;
        RECT 36.960 188.020 37.130 189.060 ;
        RECT 37.530 187.650 37.700 189.740 ;
        RECT 6.180 187.480 37.700 187.650 ;
        RECT 35.180 182.110 40.660 182.280 ;
        RECT 17.030 181.060 19.630 181.065 ;
        RECT 6.200 180.890 11.230 181.060 ;
        RECT 6.200 171.750 6.370 180.890 ;
        RECT 7.000 180.375 8.000 180.545 ;
        RECT 6.770 172.120 6.940 180.160 ;
        RECT 8.060 172.120 8.230 180.160 ;
        RECT 8.630 171.750 8.800 180.890 ;
        RECT 9.430 180.375 10.430 180.545 ;
        RECT 9.200 172.120 9.370 180.160 ;
        RECT 10.490 172.120 10.660 180.160 ;
        RECT 11.060 171.750 11.230 180.890 ;
        RECT 6.200 171.580 11.230 171.750 ;
        RECT 11.600 180.840 14.200 181.010 ;
        RECT 11.600 171.750 11.770 180.840 ;
        RECT 12.400 180.330 13.400 180.500 ;
        RECT 12.170 172.120 12.340 180.160 ;
        RECT 13.460 172.120 13.630 180.160 ;
        RECT 14.030 171.750 14.200 180.840 ;
        RECT 11.600 171.580 14.200 171.750 ;
        RECT 14.600 180.895 19.630 181.060 ;
        RECT 14.600 180.890 17.200 180.895 ;
        RECT 14.600 171.750 14.770 180.890 ;
        RECT 15.400 180.375 16.400 180.545 ;
        RECT 15.170 172.120 15.340 180.160 ;
        RECT 16.460 172.120 16.630 180.160 ;
        RECT 17.030 171.755 17.200 180.890 ;
        RECT 17.830 180.380 18.830 180.550 ;
        RECT 17.600 172.125 17.770 180.165 ;
        RECT 18.890 172.125 19.060 180.165 ;
        RECT 19.460 171.755 19.630 180.895 ;
        RECT 17.030 171.750 19.630 171.755 ;
        RECT 14.600 171.585 19.630 171.750 ;
        RECT 20.010 180.855 22.610 181.025 ;
        RECT 20.010 171.765 20.180 180.855 ;
        RECT 20.810 180.345 21.810 180.515 ;
        RECT 20.580 172.135 20.750 180.175 ;
        RECT 21.870 172.135 22.040 180.175 ;
        RECT 22.440 171.765 22.610 180.855 ;
        RECT 20.010 171.595 22.610 171.765 ;
        RECT 23.000 180.890 32.795 181.060 ;
        RECT 23.000 171.750 23.170 180.890 ;
        RECT 23.800 180.375 24.800 180.545 ;
        RECT 23.570 172.120 23.740 180.160 ;
        RECT 24.860 172.120 25.030 180.160 ;
        RECT 25.400 171.750 25.600 180.890 ;
        RECT 26.200 180.375 27.200 180.545 ;
        RECT 25.970 172.120 26.140 180.160 ;
        RECT 27.260 172.120 27.430 180.160 ;
        RECT 27.800 171.750 28.000 180.890 ;
        RECT 28.600 180.375 29.600 180.545 ;
        RECT 28.370 172.120 28.540 180.160 ;
        RECT 29.660 172.120 29.830 180.160 ;
        RECT 30.195 171.750 30.400 180.890 ;
        RECT 30.995 180.375 31.995 180.545 ;
        RECT 30.765 172.120 30.935 180.160 ;
        RECT 32.055 172.120 32.225 180.160 ;
        RECT 32.625 176.480 32.795 180.890 ;
        RECT 35.180 180.350 35.350 182.110 ;
        RECT 35.720 181.540 39.760 181.710 ;
        RECT 39.975 180.980 40.145 181.480 ;
        RECT 35.720 180.750 39.760 180.920 ;
        RECT 40.490 180.350 40.660 182.110 ;
        RECT 35.180 180.180 40.660 180.350 ;
        RECT 33.200 178.560 42.800 178.730 ;
        RECT 33.200 177.050 33.370 178.560 ;
        RECT 34.000 178.050 42.000 178.220 ;
        RECT 33.770 177.420 33.940 177.880 ;
        RECT 42.060 177.420 42.230 177.880 ;
        RECT 42.630 177.050 42.800 178.560 ;
        RECT 33.200 176.880 42.800 177.050 ;
        RECT 32.625 176.310 42.300 176.480 ;
        RECT 32.625 174.750 32.870 176.310 ;
        RECT 33.500 175.795 41.500 175.965 ;
        RECT 33.270 175.120 33.440 175.580 ;
        RECT 41.560 175.120 41.730 175.580 ;
        RECT 42.130 174.750 42.300 176.310 ;
        RECT 32.625 174.580 42.300 174.750 ;
        RECT 32.625 171.750 32.795 174.580 ;
        RECT 14.600 171.580 17.200 171.585 ;
        RECT 23.000 171.580 32.795 171.750 ;
        RECT 33.200 174.010 42.630 174.180 ;
        RECT 33.200 171.750 33.370 174.010 ;
        RECT 33.740 173.440 41.780 173.610 ;
        RECT 41.950 172.380 42.120 173.380 ;
        RECT 33.740 172.150 41.780 172.320 ;
        RECT 42.460 171.750 42.630 174.010 ;
        RECT 33.200 171.580 42.630 171.750 ;
        RECT 6.180 170.810 28.220 170.910 ;
        RECT 6.180 170.740 42.800 170.810 ;
        RECT 6.180 161.650 6.350 170.740 ;
        RECT 6.980 170.230 7.980 170.400 ;
        RECT 6.750 162.020 6.920 170.060 ;
        RECT 8.040 162.020 8.210 170.060 ;
        RECT 8.610 161.650 8.780 170.740 ;
        RECT 9.410 170.230 10.410 170.400 ;
        RECT 9.180 162.020 9.350 170.060 ;
        RECT 10.470 162.020 10.640 170.060 ;
        RECT 11.040 161.650 11.210 170.740 ;
        RECT 11.840 170.230 12.840 170.400 ;
        RECT 11.610 162.020 11.780 170.060 ;
        RECT 12.900 162.020 13.070 170.060 ;
        RECT 13.470 161.650 13.640 170.740 ;
        RECT 14.270 170.230 15.270 170.400 ;
        RECT 14.040 162.020 14.210 170.060 ;
        RECT 15.330 162.020 15.500 170.060 ;
        RECT 15.900 161.650 16.070 170.740 ;
        RECT 16.700 170.230 17.700 170.400 ;
        RECT 16.470 162.020 16.640 170.060 ;
        RECT 17.760 162.020 17.930 170.060 ;
        RECT 18.330 161.650 18.500 170.740 ;
        RECT 19.130 170.230 20.130 170.400 ;
        RECT 18.900 162.020 19.070 170.060 ;
        RECT 20.190 162.020 20.360 170.060 ;
        RECT 20.760 161.650 20.930 170.740 ;
        RECT 21.560 170.230 22.560 170.400 ;
        RECT 21.330 162.020 21.500 170.060 ;
        RECT 22.620 162.020 22.790 170.060 ;
        RECT 23.190 161.650 23.360 170.740 ;
        RECT 23.990 170.230 24.990 170.400 ;
        RECT 23.760 162.020 23.930 170.060 ;
        RECT 25.050 162.020 25.220 170.060 ;
        RECT 25.620 161.650 25.790 170.740 ;
        RECT 28.050 170.640 42.800 170.740 ;
        RECT 26.420 170.230 27.420 170.400 ;
        RECT 26.190 162.020 26.360 170.060 ;
        RECT 27.480 162.020 27.650 170.060 ;
        RECT 28.050 168.550 28.270 170.640 ;
        RECT 28.900 170.130 42.000 170.300 ;
        RECT 28.670 168.920 28.840 169.960 ;
        RECT 42.060 168.920 42.230 169.960 ;
        RECT 42.630 168.550 42.800 170.640 ;
        RECT 28.050 168.380 42.800 168.550 ;
        RECT 28.050 168.340 37.700 168.380 ;
        RECT 28.050 166.250 28.270 168.340 ;
        RECT 28.900 167.830 36.900 168.000 ;
        RECT 28.670 166.620 28.840 167.660 ;
        RECT 36.960 166.620 37.130 167.660 ;
        RECT 37.530 166.250 37.700 168.340 ;
        RECT 28.050 166.040 37.700 166.250 ;
        RECT 28.050 163.950 28.270 166.040 ;
        RECT 28.900 165.530 36.900 165.700 ;
        RECT 28.670 164.320 28.840 165.360 ;
        RECT 36.960 164.320 37.130 165.360 ;
        RECT 37.530 163.950 37.700 166.040 ;
        RECT 28.050 163.740 37.700 163.950 ;
        RECT 28.050 161.650 28.270 163.740 ;
        RECT 28.900 163.230 36.900 163.400 ;
        RECT 28.670 162.020 28.840 163.060 ;
        RECT 36.960 162.020 37.130 163.060 ;
        RECT 37.530 161.650 37.700 163.740 ;
        RECT 6.180 161.480 37.700 161.650 ;
        RECT 48.480 168.370 57.910 168.540 ;
        RECT 48.480 166.110 48.650 168.370 ;
        RECT 49.020 167.800 57.060 167.970 ;
        RECT 57.230 166.740 57.400 167.740 ;
        RECT 49.020 166.510 57.060 166.680 ;
        RECT 57.740 166.110 57.910 168.370 ;
        RECT 48.480 165.940 57.910 166.110 ;
        RECT 48.480 163.680 48.650 165.940 ;
        RECT 49.020 165.370 57.060 165.540 ;
        RECT 57.230 164.310 57.400 165.310 ;
        RECT 49.020 164.080 57.060 164.250 ;
        RECT 57.740 163.680 57.910 165.940 ;
        RECT 48.480 163.510 57.910 163.680 ;
        RECT 48.480 161.250 48.650 163.510 ;
        RECT 49.020 162.940 57.060 163.110 ;
        RECT 57.230 161.880 57.400 162.880 ;
        RECT 49.020 161.650 57.060 161.820 ;
        RECT 57.740 161.250 57.910 163.510 ;
        RECT 58.580 168.350 68.060 168.520 ;
        RECT 58.580 166.090 58.750 168.350 ;
        RECT 59.120 167.780 67.160 167.950 ;
        RECT 67.375 166.720 67.545 167.720 ;
        RECT 59.120 166.490 67.160 166.660 ;
        RECT 67.890 166.090 68.060 168.350 ;
        RECT 58.580 165.920 68.060 166.090 ;
        RECT 58.580 163.660 58.750 165.920 ;
        RECT 59.120 165.350 67.160 165.520 ;
        RECT 67.375 164.290 67.545 165.290 ;
        RECT 59.120 164.060 67.160 164.230 ;
        RECT 67.890 163.660 68.060 165.920 ;
        RECT 58.580 163.490 68.060 163.660 ;
        RECT 74.480 168.370 83.910 168.540 ;
        RECT 74.480 166.110 74.650 168.370 ;
        RECT 75.020 167.800 83.060 167.970 ;
        RECT 83.230 166.740 83.400 167.740 ;
        RECT 75.020 166.510 83.060 166.680 ;
        RECT 83.740 166.110 83.910 168.370 ;
        RECT 74.480 165.940 83.910 166.110 ;
        RECT 74.480 163.680 74.650 165.940 ;
        RECT 75.020 165.370 83.060 165.540 ;
        RECT 83.230 164.310 83.400 165.310 ;
        RECT 75.020 164.080 83.060 164.250 ;
        RECT 83.740 163.680 83.910 165.940 ;
        RECT 74.480 163.510 83.910 163.680 ;
        RECT 48.480 161.080 57.910 161.250 ;
        RECT 48.480 158.820 48.650 161.080 ;
        RECT 49.020 160.510 57.060 160.680 ;
        RECT 57.230 159.450 57.400 160.450 ;
        RECT 49.020 159.220 57.060 159.390 ;
        RECT 57.740 158.820 57.910 161.080 ;
        RECT 58.580 162.950 68.010 163.120 ;
        RECT 58.580 160.690 58.750 162.950 ;
        RECT 59.120 162.380 67.160 162.550 ;
        RECT 67.330 161.320 67.500 162.320 ;
        RECT 59.120 161.090 67.160 161.260 ;
        RECT 67.840 160.690 68.010 162.950 ;
        RECT 58.580 160.520 68.010 160.690 ;
        RECT 74.480 161.250 74.650 163.510 ;
        RECT 75.020 162.940 83.060 163.110 ;
        RECT 83.230 161.880 83.400 162.880 ;
        RECT 75.020 161.650 83.060 161.820 ;
        RECT 83.740 161.250 83.910 163.510 ;
        RECT 84.580 168.350 94.060 168.520 ;
        RECT 84.580 166.090 84.750 168.350 ;
        RECT 85.120 167.780 93.160 167.950 ;
        RECT 93.375 166.720 93.545 167.720 ;
        RECT 85.120 166.490 93.160 166.660 ;
        RECT 93.890 166.090 94.060 168.350 ;
        RECT 84.580 165.920 94.060 166.090 ;
        RECT 84.580 163.660 84.750 165.920 ;
        RECT 85.120 165.350 93.160 165.520 ;
        RECT 93.375 164.290 93.545 165.290 ;
        RECT 85.120 164.060 93.160 164.230 ;
        RECT 93.890 163.660 94.060 165.920 ;
        RECT 84.580 163.490 94.060 163.660 ;
        RECT 74.480 161.080 83.910 161.250 ;
        RECT 48.480 158.650 57.910 158.820 ;
        RECT 48.480 156.390 48.650 158.650 ;
        RECT 49.020 158.080 57.060 158.250 ;
        RECT 57.230 157.020 57.400 158.020 ;
        RECT 49.020 156.790 57.060 156.960 ;
        RECT 57.740 156.390 57.910 158.650 ;
        RECT 58.580 159.950 68.060 160.120 ;
        RECT 58.580 157.690 58.750 159.950 ;
        RECT 59.120 159.380 67.160 159.550 ;
        RECT 67.375 158.320 67.545 159.320 ;
        RECT 59.120 158.090 67.160 158.260 ;
        RECT 67.890 157.690 68.060 159.950 ;
        RECT 74.480 158.820 74.650 161.080 ;
        RECT 75.020 160.510 83.060 160.680 ;
        RECT 83.230 159.450 83.400 160.450 ;
        RECT 75.020 159.220 83.060 159.390 ;
        RECT 83.740 158.820 83.910 161.080 ;
        RECT 84.580 162.950 94.010 163.120 ;
        RECT 84.580 160.690 84.750 162.950 ;
        RECT 85.120 162.380 93.160 162.550 ;
        RECT 93.330 161.320 93.500 162.320 ;
        RECT 85.120 161.090 93.160 161.260 ;
        RECT 93.840 160.690 94.010 162.950 ;
        RECT 84.580 160.520 94.010 160.690 ;
        RECT 74.480 158.650 83.910 158.820 ;
        RECT 58.580 157.520 68.065 157.690 ;
        RECT 35.180 156.110 40.660 156.280 ;
        RECT 17.030 155.060 19.630 155.065 ;
        RECT 6.200 154.890 11.230 155.060 ;
        RECT 6.200 145.750 6.370 154.890 ;
        RECT 7.000 154.375 8.000 154.545 ;
        RECT 6.770 146.120 6.940 154.160 ;
        RECT 8.060 146.120 8.230 154.160 ;
        RECT 8.630 145.750 8.800 154.890 ;
        RECT 9.430 154.375 10.430 154.545 ;
        RECT 9.200 146.120 9.370 154.160 ;
        RECT 10.490 146.120 10.660 154.160 ;
        RECT 11.060 145.750 11.230 154.890 ;
        RECT 6.200 145.580 11.230 145.750 ;
        RECT 11.600 154.840 14.200 155.010 ;
        RECT 11.600 145.750 11.770 154.840 ;
        RECT 12.400 154.330 13.400 154.500 ;
        RECT 12.170 146.120 12.340 154.160 ;
        RECT 13.460 146.120 13.630 154.160 ;
        RECT 14.030 145.750 14.200 154.840 ;
        RECT 11.600 145.580 14.200 145.750 ;
        RECT 14.600 154.895 19.630 155.060 ;
        RECT 14.600 154.890 17.200 154.895 ;
        RECT 14.600 145.750 14.770 154.890 ;
        RECT 15.400 154.375 16.400 154.545 ;
        RECT 15.170 146.120 15.340 154.160 ;
        RECT 16.460 146.120 16.630 154.160 ;
        RECT 17.030 145.755 17.200 154.890 ;
        RECT 17.830 154.380 18.830 154.550 ;
        RECT 17.600 146.125 17.770 154.165 ;
        RECT 18.890 146.125 19.060 154.165 ;
        RECT 19.460 145.755 19.630 154.895 ;
        RECT 17.030 145.750 19.630 145.755 ;
        RECT 14.600 145.585 19.630 145.750 ;
        RECT 20.010 154.855 22.610 155.025 ;
        RECT 20.010 145.765 20.180 154.855 ;
        RECT 20.810 154.345 21.810 154.515 ;
        RECT 20.580 146.135 20.750 154.175 ;
        RECT 21.870 146.135 22.040 154.175 ;
        RECT 22.440 145.765 22.610 154.855 ;
        RECT 20.010 145.595 22.610 145.765 ;
        RECT 23.000 154.890 32.795 155.060 ;
        RECT 23.000 145.750 23.170 154.890 ;
        RECT 23.800 154.375 24.800 154.545 ;
        RECT 23.570 146.120 23.740 154.160 ;
        RECT 24.860 146.120 25.030 154.160 ;
        RECT 25.400 145.750 25.600 154.890 ;
        RECT 26.200 154.375 27.200 154.545 ;
        RECT 25.970 146.120 26.140 154.160 ;
        RECT 27.260 146.120 27.430 154.160 ;
        RECT 27.800 145.750 28.000 154.890 ;
        RECT 28.600 154.375 29.600 154.545 ;
        RECT 28.370 146.120 28.540 154.160 ;
        RECT 29.660 146.120 29.830 154.160 ;
        RECT 30.195 145.750 30.400 154.890 ;
        RECT 30.995 154.375 31.995 154.545 ;
        RECT 30.765 146.120 30.935 154.160 ;
        RECT 32.055 146.120 32.225 154.160 ;
        RECT 32.625 150.480 32.795 154.890 ;
        RECT 35.180 154.350 35.350 156.110 ;
        RECT 35.720 155.540 39.760 155.710 ;
        RECT 39.975 154.980 40.145 155.480 ;
        RECT 35.720 154.750 39.760 154.920 ;
        RECT 40.490 154.350 40.660 156.110 ;
        RECT 35.180 154.180 40.660 154.350 ;
        RECT 48.480 156.220 57.910 156.390 ;
        RECT 48.480 153.960 48.650 156.220 ;
        RECT 49.020 155.650 57.060 155.820 ;
        RECT 57.230 154.590 57.400 155.590 ;
        RECT 49.020 154.360 57.060 154.530 ;
        RECT 57.740 153.960 57.910 156.220 ;
        RECT 58.585 155.260 58.755 157.520 ;
        RECT 59.125 156.950 67.165 157.120 ;
        RECT 67.380 155.890 67.550 156.890 ;
        RECT 59.125 155.660 67.165 155.830 ;
        RECT 67.895 155.260 68.065 157.520 ;
        RECT 58.585 155.090 68.065 155.260 ;
        RECT 74.480 156.390 74.650 158.650 ;
        RECT 75.020 158.080 83.060 158.250 ;
        RECT 83.230 157.020 83.400 158.020 ;
        RECT 75.020 156.790 83.060 156.960 ;
        RECT 83.740 156.390 83.910 158.650 ;
        RECT 84.580 159.950 94.060 160.120 ;
        RECT 84.580 157.690 84.750 159.950 ;
        RECT 85.120 159.380 93.160 159.550 ;
        RECT 93.375 158.320 93.545 159.320 ;
        RECT 85.120 158.090 93.160 158.260 ;
        RECT 93.890 157.690 94.060 159.950 ;
        RECT 84.580 157.520 94.065 157.690 ;
        RECT 74.480 156.220 83.910 156.390 ;
        RECT 48.480 153.790 57.910 153.960 ;
        RECT 33.200 152.560 42.800 152.730 ;
        RECT 33.200 151.050 33.370 152.560 ;
        RECT 34.000 152.050 42.000 152.220 ;
        RECT 33.770 151.420 33.940 151.880 ;
        RECT 42.060 151.420 42.230 151.880 ;
        RECT 42.630 151.050 42.800 152.560 ;
        RECT 33.200 150.880 42.800 151.050 ;
        RECT 48.480 151.530 48.650 153.790 ;
        RECT 49.020 153.220 57.060 153.390 ;
        RECT 57.230 152.160 57.400 153.160 ;
        RECT 49.020 151.930 57.060 152.100 ;
        RECT 57.740 151.530 57.910 153.790 ;
        RECT 58.595 154.540 68.025 154.710 ;
        RECT 58.595 152.280 58.765 154.540 ;
        RECT 59.135 153.970 67.175 154.140 ;
        RECT 67.345 152.910 67.515 153.910 ;
        RECT 59.135 152.680 67.175 152.850 ;
        RECT 67.855 152.280 68.025 154.540 ;
        RECT 58.595 152.110 68.025 152.280 ;
        RECT 74.480 153.960 74.650 156.220 ;
        RECT 75.020 155.650 83.060 155.820 ;
        RECT 83.230 154.590 83.400 155.590 ;
        RECT 75.020 154.360 83.060 154.530 ;
        RECT 83.740 153.960 83.910 156.220 ;
        RECT 84.585 155.260 84.755 157.520 ;
        RECT 85.125 156.950 93.165 157.120 ;
        RECT 93.380 155.890 93.550 156.890 ;
        RECT 85.125 155.660 93.165 155.830 ;
        RECT 93.895 155.260 94.065 157.520 ;
        RECT 84.585 155.090 94.065 155.260 ;
        RECT 74.480 153.790 83.910 153.960 ;
        RECT 48.480 151.360 57.910 151.530 ;
        RECT 32.625 150.310 42.300 150.480 ;
        RECT 32.625 148.750 32.870 150.310 ;
        RECT 33.500 149.795 41.500 149.965 ;
        RECT 33.270 149.120 33.440 149.580 ;
        RECT 41.560 149.120 41.730 149.580 ;
        RECT 42.130 148.750 42.300 150.310 ;
        RECT 32.625 148.580 42.300 148.750 ;
        RECT 48.480 149.100 48.650 151.360 ;
        RECT 49.020 150.790 57.060 150.960 ;
        RECT 57.230 149.730 57.400 150.730 ;
        RECT 49.020 149.500 57.060 149.670 ;
        RECT 57.740 149.100 57.910 151.360 ;
        RECT 48.480 148.930 57.910 149.100 ;
        RECT 32.625 145.750 32.795 148.580 ;
        RECT 14.600 145.580 17.200 145.585 ;
        RECT 23.000 145.580 32.795 145.750 ;
        RECT 33.200 148.010 42.630 148.180 ;
        RECT 33.200 145.750 33.370 148.010 ;
        RECT 33.740 147.440 41.780 147.610 ;
        RECT 41.950 146.380 42.120 147.380 ;
        RECT 33.740 146.150 41.780 146.320 ;
        RECT 42.460 145.750 42.630 148.010 ;
        RECT 33.200 145.580 42.630 145.750 ;
        RECT 48.480 146.670 48.650 148.930 ;
        RECT 49.020 148.360 57.060 148.530 ;
        RECT 57.230 147.300 57.400 148.300 ;
        RECT 49.020 147.070 57.060 147.240 ;
        RECT 57.740 146.670 57.910 148.930 ;
        RECT 48.480 146.500 57.910 146.670 ;
        RECT 58.580 151.550 68.060 151.720 ;
        RECT 58.580 149.320 58.750 151.550 ;
        RECT 59.120 150.980 67.160 151.150 ;
        RECT 67.375 149.920 67.545 150.920 ;
        RECT 59.120 149.690 67.160 149.860 ;
        RECT 67.890 149.320 68.060 151.550 ;
        RECT 58.580 149.120 68.060 149.320 ;
        RECT 58.580 146.920 58.750 149.120 ;
        RECT 59.120 148.580 67.160 148.750 ;
        RECT 67.375 147.520 67.545 148.520 ;
        RECT 59.120 147.290 67.160 147.460 ;
        RECT 67.890 146.920 68.060 149.120 ;
        RECT 58.580 146.720 68.060 146.920 ;
        RECT 48.480 146.450 57.810 146.500 ;
        RECT 6.180 144.810 28.220 144.910 ;
        RECT 6.180 144.740 42.800 144.810 ;
        RECT 6.180 135.650 6.350 144.740 ;
        RECT 6.980 144.230 7.980 144.400 ;
        RECT 6.750 136.020 6.920 144.060 ;
        RECT 8.040 136.020 8.210 144.060 ;
        RECT 8.610 135.650 8.780 144.740 ;
        RECT 9.410 144.230 10.410 144.400 ;
        RECT 9.180 136.020 9.350 144.060 ;
        RECT 10.470 136.020 10.640 144.060 ;
        RECT 11.040 135.650 11.210 144.740 ;
        RECT 11.840 144.230 12.840 144.400 ;
        RECT 11.610 136.020 11.780 144.060 ;
        RECT 12.900 136.020 13.070 144.060 ;
        RECT 13.470 135.650 13.640 144.740 ;
        RECT 14.270 144.230 15.270 144.400 ;
        RECT 14.040 136.020 14.210 144.060 ;
        RECT 15.330 136.020 15.500 144.060 ;
        RECT 15.900 135.650 16.070 144.740 ;
        RECT 16.700 144.230 17.700 144.400 ;
        RECT 16.470 136.020 16.640 144.060 ;
        RECT 17.760 136.020 17.930 144.060 ;
        RECT 18.330 135.650 18.500 144.740 ;
        RECT 19.130 144.230 20.130 144.400 ;
        RECT 18.900 136.020 19.070 144.060 ;
        RECT 20.190 136.020 20.360 144.060 ;
        RECT 20.760 135.650 20.930 144.740 ;
        RECT 21.560 144.230 22.560 144.400 ;
        RECT 21.330 136.020 21.500 144.060 ;
        RECT 22.620 136.020 22.790 144.060 ;
        RECT 23.190 135.650 23.360 144.740 ;
        RECT 23.990 144.230 24.990 144.400 ;
        RECT 23.760 136.020 23.930 144.060 ;
        RECT 25.050 136.020 25.220 144.060 ;
        RECT 25.620 135.650 25.790 144.740 ;
        RECT 28.050 144.640 42.800 144.740 ;
        RECT 26.420 144.230 27.420 144.400 ;
        RECT 26.190 136.020 26.360 144.060 ;
        RECT 27.480 136.020 27.650 144.060 ;
        RECT 28.050 142.550 28.270 144.640 ;
        RECT 28.900 144.130 42.000 144.300 ;
        RECT 28.670 142.920 28.840 143.960 ;
        RECT 42.060 142.920 42.230 143.960 ;
        RECT 42.630 142.550 42.800 144.640 ;
        RECT 28.050 142.380 42.800 142.550 ;
        RECT 28.050 142.340 37.700 142.380 ;
        RECT 28.050 140.250 28.270 142.340 ;
        RECT 28.900 141.830 36.900 142.000 ;
        RECT 28.670 140.620 28.840 141.660 ;
        RECT 36.960 140.620 37.130 141.660 ;
        RECT 37.530 140.250 37.700 142.340 ;
        RECT 28.050 140.040 37.700 140.250 ;
        RECT 28.050 137.950 28.270 140.040 ;
        RECT 28.900 139.530 36.900 139.700 ;
        RECT 28.670 138.320 28.840 139.360 ;
        RECT 36.960 138.320 37.130 139.360 ;
        RECT 37.530 137.950 37.700 140.040 ;
        RECT 28.050 137.740 37.700 137.950 ;
        RECT 28.050 135.650 28.270 137.740 ;
        RECT 28.900 137.230 36.900 137.400 ;
        RECT 28.670 136.020 28.840 137.060 ;
        RECT 36.960 136.020 37.130 137.060 ;
        RECT 37.530 135.650 37.700 137.740 ;
        RECT 48.480 137.190 48.650 146.450 ;
        RECT 49.020 145.880 50.060 146.050 ;
        RECT 50.230 137.820 50.400 145.820 ;
        RECT 49.020 137.590 50.060 137.760 ;
        RECT 50.740 137.190 50.950 146.450 ;
        RECT 51.320 145.880 52.360 146.050 ;
        RECT 52.530 137.820 52.700 145.820 ;
        RECT 51.320 137.590 52.360 137.760 ;
        RECT 53.040 137.190 53.250 146.450 ;
        RECT 53.620 145.880 54.660 146.050 ;
        RECT 54.830 137.820 55.000 145.820 ;
        RECT 53.620 137.590 54.660 137.760 ;
        RECT 55.340 137.190 55.550 146.450 ;
        RECT 55.920 145.880 56.960 146.050 ;
        RECT 48.480 137.020 55.550 137.190 ;
        RECT 6.180 135.480 37.700 135.650 ;
        RECT 55.380 132.090 55.550 137.020 ;
        RECT 57.130 132.720 57.300 145.820 ;
        RECT 55.920 132.490 56.960 132.660 ;
        RECT 57.640 132.090 57.810 146.450 ;
        RECT 58.580 144.525 58.750 146.720 ;
        RECT 59.120 146.180 67.160 146.350 ;
        RECT 67.375 145.120 67.545 146.120 ;
        RECT 59.120 144.890 67.160 145.060 ;
        RECT 67.890 144.525 68.060 146.720 ;
        RECT 58.580 144.320 68.060 144.525 ;
        RECT 58.580 142.095 58.750 144.320 ;
        RECT 59.120 143.785 67.160 143.955 ;
        RECT 67.375 142.725 67.545 143.725 ;
        RECT 59.120 142.495 67.160 142.665 ;
        RECT 67.890 142.095 68.060 144.320 ;
        RECT 58.580 141.925 68.060 142.095 ;
        RECT 74.480 151.530 74.650 153.790 ;
        RECT 75.020 153.220 83.060 153.390 ;
        RECT 83.230 152.160 83.400 153.160 ;
        RECT 75.020 151.930 83.060 152.100 ;
        RECT 83.740 151.530 83.910 153.790 ;
        RECT 84.595 154.540 94.025 154.710 ;
        RECT 84.595 152.280 84.765 154.540 ;
        RECT 85.135 153.970 93.175 154.140 ;
        RECT 93.345 152.910 93.515 153.910 ;
        RECT 85.135 152.680 93.175 152.850 ;
        RECT 93.855 152.280 94.025 154.540 ;
        RECT 84.595 152.110 94.025 152.280 ;
        RECT 74.480 151.360 83.910 151.530 ;
        RECT 74.480 149.100 74.650 151.360 ;
        RECT 75.020 150.790 83.060 150.960 ;
        RECT 83.230 149.730 83.400 150.730 ;
        RECT 75.020 149.500 83.060 149.670 ;
        RECT 83.740 149.100 83.910 151.360 ;
        RECT 74.480 148.930 83.910 149.100 ;
        RECT 74.480 146.670 74.650 148.930 ;
        RECT 75.020 148.360 83.060 148.530 ;
        RECT 83.230 147.300 83.400 148.300 ;
        RECT 75.020 147.070 83.060 147.240 ;
        RECT 83.740 146.670 83.910 148.930 ;
        RECT 74.480 146.500 83.910 146.670 ;
        RECT 84.580 151.550 94.060 151.720 ;
        RECT 84.580 149.320 84.750 151.550 ;
        RECT 85.120 150.980 93.160 151.150 ;
        RECT 93.375 149.920 93.545 150.920 ;
        RECT 85.120 149.690 93.160 149.860 ;
        RECT 93.890 149.320 94.060 151.550 ;
        RECT 84.580 149.120 94.060 149.320 ;
        RECT 84.580 146.920 84.750 149.120 ;
        RECT 85.120 148.580 93.160 148.750 ;
        RECT 93.375 147.520 93.545 148.520 ;
        RECT 85.120 147.290 93.160 147.460 ;
        RECT 93.890 146.920 94.060 149.120 ;
        RECT 84.580 146.720 94.060 146.920 ;
        RECT 74.480 146.450 83.810 146.500 ;
        RECT 61.580 141.850 63.480 141.925 ;
        RECT 58.580 141.350 61.180 141.520 ;
        RECT 58.580 132.260 58.750 141.350 ;
        RECT 59.150 132.940 59.320 140.980 ;
        RECT 60.440 132.940 60.610 140.980 ;
        RECT 59.380 132.600 60.380 132.770 ;
        RECT 61.010 132.260 61.180 141.350 ;
        RECT 61.580 132.590 61.750 141.850 ;
        RECT 62.120 141.280 62.580 141.450 ;
        RECT 62.795 133.220 62.965 141.220 ;
        RECT 62.120 132.990 62.580 133.160 ;
        RECT 63.310 132.590 63.480 141.850 ;
        RECT 61.580 132.420 63.480 132.590 ;
        RECT 63.880 141.350 65.730 141.520 ;
        RECT 58.580 132.090 61.180 132.260 ;
        RECT 63.880 132.090 64.050 141.350 ;
        RECT 64.420 140.780 64.880 140.950 ;
        RECT 65.050 132.720 65.220 140.720 ;
        RECT 64.420 132.490 64.880 132.660 ;
        RECT 65.560 132.090 65.730 141.350 ;
        RECT 67.180 139.490 69.280 139.660 ;
        RECT 67.180 134.350 67.350 139.490 ;
        RECT 67.750 135.080 67.920 139.120 ;
        RECT 68.540 135.080 68.710 139.120 ;
        RECT 67.980 134.695 68.480 134.865 ;
        RECT 69.110 134.350 69.280 139.490 ;
        RECT 74.480 137.190 74.650 146.450 ;
        RECT 75.020 145.880 76.060 146.050 ;
        RECT 76.230 137.820 76.400 145.820 ;
        RECT 75.020 137.590 76.060 137.760 ;
        RECT 76.740 137.190 76.950 146.450 ;
        RECT 77.320 145.880 78.360 146.050 ;
        RECT 78.530 137.820 78.700 145.820 ;
        RECT 77.320 137.590 78.360 137.760 ;
        RECT 79.040 137.190 79.250 146.450 ;
        RECT 79.620 145.880 80.660 146.050 ;
        RECT 80.830 137.820 81.000 145.820 ;
        RECT 79.620 137.590 80.660 137.760 ;
        RECT 81.340 137.190 81.550 146.450 ;
        RECT 81.920 145.880 82.960 146.050 ;
        RECT 74.480 137.020 81.550 137.190 ;
        RECT 67.180 134.180 69.280 134.350 ;
        RECT 55.380 131.920 57.810 132.090 ;
        RECT 63.880 131.920 65.730 132.090 ;
        RECT 81.380 132.090 81.550 137.020 ;
        RECT 83.130 132.720 83.300 145.820 ;
        RECT 81.920 132.490 82.960 132.660 ;
        RECT 83.640 132.090 83.810 146.450 ;
        RECT 84.580 144.525 84.750 146.720 ;
        RECT 85.120 146.180 93.160 146.350 ;
        RECT 93.375 145.120 93.545 146.120 ;
        RECT 85.120 144.890 93.160 145.060 ;
        RECT 93.890 144.525 94.060 146.720 ;
        RECT 84.580 144.320 94.060 144.525 ;
        RECT 84.580 142.095 84.750 144.320 ;
        RECT 85.120 143.785 93.160 143.955 ;
        RECT 93.375 142.725 93.545 143.725 ;
        RECT 85.120 142.495 93.160 142.665 ;
        RECT 93.890 142.095 94.060 144.320 ;
        RECT 84.580 141.925 94.060 142.095 ;
        RECT 87.580 141.850 89.480 141.925 ;
        RECT 84.580 141.350 87.180 141.520 ;
        RECT 84.580 132.260 84.750 141.350 ;
        RECT 85.150 132.940 85.320 140.980 ;
        RECT 86.440 132.940 86.610 140.980 ;
        RECT 85.380 132.600 86.380 132.770 ;
        RECT 87.010 132.260 87.180 141.350 ;
        RECT 87.580 132.590 87.750 141.850 ;
        RECT 88.120 141.280 88.580 141.450 ;
        RECT 88.795 133.220 88.965 141.220 ;
        RECT 88.120 132.990 88.580 133.160 ;
        RECT 89.310 132.590 89.480 141.850 ;
        RECT 87.580 132.420 89.480 132.590 ;
        RECT 89.880 141.350 91.730 141.520 ;
        RECT 84.580 132.090 87.180 132.260 ;
        RECT 89.880 132.090 90.050 141.350 ;
        RECT 90.420 140.780 90.880 140.950 ;
        RECT 91.050 132.720 91.220 140.720 ;
        RECT 90.420 132.490 90.880 132.660 ;
        RECT 91.560 132.090 91.730 141.350 ;
        RECT 93.180 139.490 95.280 139.660 ;
        RECT 93.180 134.350 93.350 139.490 ;
        RECT 93.750 135.080 93.920 139.120 ;
        RECT 94.540 135.080 94.710 139.120 ;
        RECT 93.980 134.695 94.480 134.865 ;
        RECT 95.110 134.350 95.280 139.490 ;
        RECT 93.180 134.180 95.280 134.350 ;
        RECT 81.380 131.920 83.810 132.090 ;
        RECT 89.880 131.920 91.730 132.090 ;
        RECT 35.180 130.110 40.660 130.280 ;
        RECT 17.030 129.060 19.630 129.065 ;
        RECT 6.200 128.890 11.230 129.060 ;
        RECT 6.200 119.750 6.370 128.890 ;
        RECT 7.000 128.375 8.000 128.545 ;
        RECT 6.770 120.120 6.940 128.160 ;
        RECT 8.060 120.120 8.230 128.160 ;
        RECT 8.630 119.750 8.800 128.890 ;
        RECT 9.430 128.375 10.430 128.545 ;
        RECT 9.200 120.120 9.370 128.160 ;
        RECT 10.490 120.120 10.660 128.160 ;
        RECT 11.060 119.750 11.230 128.890 ;
        RECT 6.200 119.580 11.230 119.750 ;
        RECT 11.600 128.840 14.200 129.010 ;
        RECT 11.600 119.750 11.770 128.840 ;
        RECT 12.400 128.330 13.400 128.500 ;
        RECT 12.170 120.120 12.340 128.160 ;
        RECT 13.460 120.120 13.630 128.160 ;
        RECT 14.030 119.750 14.200 128.840 ;
        RECT 11.600 119.580 14.200 119.750 ;
        RECT 14.600 128.895 19.630 129.060 ;
        RECT 14.600 128.890 17.200 128.895 ;
        RECT 14.600 119.750 14.770 128.890 ;
        RECT 15.400 128.375 16.400 128.545 ;
        RECT 15.170 120.120 15.340 128.160 ;
        RECT 16.460 120.120 16.630 128.160 ;
        RECT 17.030 119.755 17.200 128.890 ;
        RECT 17.830 128.380 18.830 128.550 ;
        RECT 17.600 120.125 17.770 128.165 ;
        RECT 18.890 120.125 19.060 128.165 ;
        RECT 19.460 119.755 19.630 128.895 ;
        RECT 17.030 119.750 19.630 119.755 ;
        RECT 14.600 119.585 19.630 119.750 ;
        RECT 20.010 128.855 22.610 129.025 ;
        RECT 20.010 119.765 20.180 128.855 ;
        RECT 20.810 128.345 21.810 128.515 ;
        RECT 20.580 120.135 20.750 128.175 ;
        RECT 21.870 120.135 22.040 128.175 ;
        RECT 22.440 119.765 22.610 128.855 ;
        RECT 20.010 119.595 22.610 119.765 ;
        RECT 23.000 128.890 32.795 129.060 ;
        RECT 23.000 119.750 23.170 128.890 ;
        RECT 23.800 128.375 24.800 128.545 ;
        RECT 23.570 120.120 23.740 128.160 ;
        RECT 24.860 120.120 25.030 128.160 ;
        RECT 25.400 119.750 25.600 128.890 ;
        RECT 26.200 128.375 27.200 128.545 ;
        RECT 25.970 120.120 26.140 128.160 ;
        RECT 27.260 120.120 27.430 128.160 ;
        RECT 27.800 119.750 28.000 128.890 ;
        RECT 28.600 128.375 29.600 128.545 ;
        RECT 28.370 120.120 28.540 128.160 ;
        RECT 29.660 120.120 29.830 128.160 ;
        RECT 30.195 119.750 30.400 128.890 ;
        RECT 30.995 128.375 31.995 128.545 ;
        RECT 30.765 120.120 30.935 128.160 ;
        RECT 32.055 120.120 32.225 128.160 ;
        RECT 32.625 124.480 32.795 128.890 ;
        RECT 35.180 128.350 35.350 130.110 ;
        RECT 35.720 129.540 39.760 129.710 ;
        RECT 39.975 128.980 40.145 129.480 ;
        RECT 35.720 128.750 39.760 128.920 ;
        RECT 40.490 128.350 40.660 130.110 ;
        RECT 35.180 128.180 40.660 128.350 ;
        RECT 33.200 126.560 42.800 126.730 ;
        RECT 33.200 125.050 33.370 126.560 ;
        RECT 34.000 126.050 42.000 126.220 ;
        RECT 33.770 125.420 33.940 125.880 ;
        RECT 42.060 125.420 42.230 125.880 ;
        RECT 42.630 125.050 42.800 126.560 ;
        RECT 33.200 124.880 42.800 125.050 ;
        RECT 48.480 126.370 57.910 126.540 ;
        RECT 32.625 124.310 42.300 124.480 ;
        RECT 32.625 122.750 32.870 124.310 ;
        RECT 33.500 123.795 41.500 123.965 ;
        RECT 33.270 123.120 33.440 123.580 ;
        RECT 41.560 123.120 41.730 123.580 ;
        RECT 42.130 122.750 42.300 124.310 ;
        RECT 32.625 122.580 42.300 122.750 ;
        RECT 48.480 124.110 48.650 126.370 ;
        RECT 49.020 125.800 57.060 125.970 ;
        RECT 57.230 124.740 57.400 125.740 ;
        RECT 49.020 124.510 57.060 124.680 ;
        RECT 57.740 124.110 57.910 126.370 ;
        RECT 48.480 123.940 57.910 124.110 ;
        RECT 32.625 119.750 32.795 122.580 ;
        RECT 14.600 119.580 17.200 119.585 ;
        RECT 23.000 119.580 32.795 119.750 ;
        RECT 33.200 122.010 42.630 122.180 ;
        RECT 33.200 119.750 33.370 122.010 ;
        RECT 33.740 121.440 41.780 121.610 ;
        RECT 41.950 120.380 42.120 121.380 ;
        RECT 33.740 120.150 41.780 120.320 ;
        RECT 42.460 119.750 42.630 122.010 ;
        RECT 33.200 119.580 42.630 119.750 ;
        RECT 48.480 121.680 48.650 123.940 ;
        RECT 49.020 123.370 57.060 123.540 ;
        RECT 57.230 122.310 57.400 123.310 ;
        RECT 49.020 122.080 57.060 122.250 ;
        RECT 57.740 121.680 57.910 123.940 ;
        RECT 48.480 121.510 57.910 121.680 ;
        RECT 48.480 119.250 48.650 121.510 ;
        RECT 49.020 120.940 57.060 121.110 ;
        RECT 57.230 119.880 57.400 120.880 ;
        RECT 49.020 119.650 57.060 119.820 ;
        RECT 57.740 119.250 57.910 121.510 ;
        RECT 58.580 126.350 68.060 126.520 ;
        RECT 58.580 124.090 58.750 126.350 ;
        RECT 59.120 125.780 67.160 125.950 ;
        RECT 67.375 124.720 67.545 125.720 ;
        RECT 59.120 124.490 67.160 124.660 ;
        RECT 67.890 124.090 68.060 126.350 ;
        RECT 58.580 123.920 68.060 124.090 ;
        RECT 58.580 121.660 58.750 123.920 ;
        RECT 59.120 123.350 67.160 123.520 ;
        RECT 67.375 122.290 67.545 123.290 ;
        RECT 59.120 122.060 67.160 122.230 ;
        RECT 67.890 121.660 68.060 123.920 ;
        RECT 58.580 121.490 68.060 121.660 ;
        RECT 74.480 126.370 83.910 126.540 ;
        RECT 74.480 124.110 74.650 126.370 ;
        RECT 75.020 125.800 83.060 125.970 ;
        RECT 83.230 124.740 83.400 125.740 ;
        RECT 75.020 124.510 83.060 124.680 ;
        RECT 83.740 124.110 83.910 126.370 ;
        RECT 74.480 123.940 83.910 124.110 ;
        RECT 74.480 121.680 74.650 123.940 ;
        RECT 75.020 123.370 83.060 123.540 ;
        RECT 83.230 122.310 83.400 123.310 ;
        RECT 75.020 122.080 83.060 122.250 ;
        RECT 83.740 121.680 83.910 123.940 ;
        RECT 74.480 121.510 83.910 121.680 ;
        RECT 48.480 119.080 57.910 119.250 ;
        RECT 6.180 118.810 28.220 118.910 ;
        RECT 6.180 118.740 42.800 118.810 ;
        RECT 6.180 109.650 6.350 118.740 ;
        RECT 6.980 118.230 7.980 118.400 ;
        RECT 6.750 110.020 6.920 118.060 ;
        RECT 8.040 110.020 8.210 118.060 ;
        RECT 8.610 109.650 8.780 118.740 ;
        RECT 9.410 118.230 10.410 118.400 ;
        RECT 9.180 110.020 9.350 118.060 ;
        RECT 10.470 110.020 10.640 118.060 ;
        RECT 11.040 109.650 11.210 118.740 ;
        RECT 11.840 118.230 12.840 118.400 ;
        RECT 11.610 110.020 11.780 118.060 ;
        RECT 12.900 110.020 13.070 118.060 ;
        RECT 13.470 109.650 13.640 118.740 ;
        RECT 14.270 118.230 15.270 118.400 ;
        RECT 14.040 110.020 14.210 118.060 ;
        RECT 15.330 110.020 15.500 118.060 ;
        RECT 15.900 109.650 16.070 118.740 ;
        RECT 16.700 118.230 17.700 118.400 ;
        RECT 16.470 110.020 16.640 118.060 ;
        RECT 17.760 110.020 17.930 118.060 ;
        RECT 18.330 109.650 18.500 118.740 ;
        RECT 19.130 118.230 20.130 118.400 ;
        RECT 18.900 110.020 19.070 118.060 ;
        RECT 20.190 110.020 20.360 118.060 ;
        RECT 20.760 109.650 20.930 118.740 ;
        RECT 21.560 118.230 22.560 118.400 ;
        RECT 21.330 110.020 21.500 118.060 ;
        RECT 22.620 110.020 22.790 118.060 ;
        RECT 23.190 109.650 23.360 118.740 ;
        RECT 23.990 118.230 24.990 118.400 ;
        RECT 23.760 110.020 23.930 118.060 ;
        RECT 25.050 110.020 25.220 118.060 ;
        RECT 25.620 109.650 25.790 118.740 ;
        RECT 28.050 118.640 42.800 118.740 ;
        RECT 26.420 118.230 27.420 118.400 ;
        RECT 26.190 110.020 26.360 118.060 ;
        RECT 27.480 110.020 27.650 118.060 ;
        RECT 28.050 116.550 28.270 118.640 ;
        RECT 28.900 118.130 42.000 118.300 ;
        RECT 28.670 116.920 28.840 117.960 ;
        RECT 42.060 116.920 42.230 117.960 ;
        RECT 42.630 116.550 42.800 118.640 ;
        RECT 28.050 116.380 42.800 116.550 ;
        RECT 48.480 116.820 48.650 119.080 ;
        RECT 49.020 118.510 57.060 118.680 ;
        RECT 57.230 117.450 57.400 118.450 ;
        RECT 49.020 117.220 57.060 117.390 ;
        RECT 57.740 116.820 57.910 119.080 ;
        RECT 58.580 120.950 68.010 121.120 ;
        RECT 58.580 118.690 58.750 120.950 ;
        RECT 59.120 120.380 67.160 120.550 ;
        RECT 67.330 119.320 67.500 120.320 ;
        RECT 59.120 119.090 67.160 119.260 ;
        RECT 67.840 118.690 68.010 120.950 ;
        RECT 58.580 118.520 68.010 118.690 ;
        RECT 74.480 119.250 74.650 121.510 ;
        RECT 75.020 120.940 83.060 121.110 ;
        RECT 83.230 119.880 83.400 120.880 ;
        RECT 75.020 119.650 83.060 119.820 ;
        RECT 83.740 119.250 83.910 121.510 ;
        RECT 84.580 126.350 94.060 126.520 ;
        RECT 84.580 124.090 84.750 126.350 ;
        RECT 85.120 125.780 93.160 125.950 ;
        RECT 93.375 124.720 93.545 125.720 ;
        RECT 85.120 124.490 93.160 124.660 ;
        RECT 93.890 124.090 94.060 126.350 ;
        RECT 84.580 123.920 94.060 124.090 ;
        RECT 84.580 121.660 84.750 123.920 ;
        RECT 85.120 123.350 93.160 123.520 ;
        RECT 93.375 122.290 93.545 123.290 ;
        RECT 85.120 122.060 93.160 122.230 ;
        RECT 93.890 121.660 94.060 123.920 ;
        RECT 84.580 121.490 94.060 121.660 ;
        RECT 74.480 119.080 83.910 119.250 ;
        RECT 48.480 116.650 57.910 116.820 ;
        RECT 28.050 116.340 37.700 116.380 ;
        RECT 28.050 114.250 28.270 116.340 ;
        RECT 28.900 115.830 36.900 116.000 ;
        RECT 28.670 114.620 28.840 115.660 ;
        RECT 36.960 114.620 37.130 115.660 ;
        RECT 37.530 114.250 37.700 116.340 ;
        RECT 28.050 114.040 37.700 114.250 ;
        RECT 28.050 111.950 28.270 114.040 ;
        RECT 28.900 113.530 36.900 113.700 ;
        RECT 28.670 112.320 28.840 113.360 ;
        RECT 36.960 112.320 37.130 113.360 ;
        RECT 37.530 111.950 37.700 114.040 ;
        RECT 28.050 111.740 37.700 111.950 ;
        RECT 28.050 109.650 28.270 111.740 ;
        RECT 28.900 111.230 36.900 111.400 ;
        RECT 28.670 110.020 28.840 111.060 ;
        RECT 36.960 110.020 37.130 111.060 ;
        RECT 37.530 109.650 37.700 111.740 ;
        RECT 6.180 109.480 37.700 109.650 ;
        RECT 48.480 114.390 48.650 116.650 ;
        RECT 49.020 116.080 57.060 116.250 ;
        RECT 57.230 115.020 57.400 116.020 ;
        RECT 49.020 114.790 57.060 114.960 ;
        RECT 57.740 114.390 57.910 116.650 ;
        RECT 58.580 117.950 68.060 118.120 ;
        RECT 58.580 115.690 58.750 117.950 ;
        RECT 59.120 117.380 67.160 117.550 ;
        RECT 67.375 116.320 67.545 117.320 ;
        RECT 59.120 116.090 67.160 116.260 ;
        RECT 67.890 115.690 68.060 117.950 ;
        RECT 74.480 116.820 74.650 119.080 ;
        RECT 75.020 118.510 83.060 118.680 ;
        RECT 83.230 117.450 83.400 118.450 ;
        RECT 75.020 117.220 83.060 117.390 ;
        RECT 83.740 116.820 83.910 119.080 ;
        RECT 84.580 120.950 94.010 121.120 ;
        RECT 84.580 118.690 84.750 120.950 ;
        RECT 85.120 120.380 93.160 120.550 ;
        RECT 93.330 119.320 93.500 120.320 ;
        RECT 85.120 119.090 93.160 119.260 ;
        RECT 93.840 118.690 94.010 120.950 ;
        RECT 84.580 118.520 94.010 118.690 ;
        RECT 74.480 116.650 83.910 116.820 ;
        RECT 58.580 115.520 68.065 115.690 ;
        RECT 48.480 114.220 57.910 114.390 ;
        RECT 48.480 111.960 48.650 114.220 ;
        RECT 49.020 113.650 57.060 113.820 ;
        RECT 57.230 112.590 57.400 113.590 ;
        RECT 49.020 112.360 57.060 112.530 ;
        RECT 57.740 111.960 57.910 114.220 ;
        RECT 58.585 113.260 58.755 115.520 ;
        RECT 59.125 114.950 67.165 115.120 ;
        RECT 67.380 113.890 67.550 114.890 ;
        RECT 59.125 113.660 67.165 113.830 ;
        RECT 67.895 113.260 68.065 115.520 ;
        RECT 58.585 113.090 68.065 113.260 ;
        RECT 74.480 114.390 74.650 116.650 ;
        RECT 75.020 116.080 83.060 116.250 ;
        RECT 83.230 115.020 83.400 116.020 ;
        RECT 75.020 114.790 83.060 114.960 ;
        RECT 83.740 114.390 83.910 116.650 ;
        RECT 84.580 117.950 94.060 118.120 ;
        RECT 84.580 115.690 84.750 117.950 ;
        RECT 85.120 117.380 93.160 117.550 ;
        RECT 93.375 116.320 93.545 117.320 ;
        RECT 85.120 116.090 93.160 116.260 ;
        RECT 93.890 115.690 94.060 117.950 ;
        RECT 84.580 115.520 94.065 115.690 ;
        RECT 74.480 114.220 83.910 114.390 ;
        RECT 48.480 111.790 57.910 111.960 ;
        RECT 48.480 109.530 48.650 111.790 ;
        RECT 49.020 111.220 57.060 111.390 ;
        RECT 57.230 110.160 57.400 111.160 ;
        RECT 49.020 109.930 57.060 110.100 ;
        RECT 57.740 109.530 57.910 111.790 ;
        RECT 58.595 112.540 68.025 112.710 ;
        RECT 58.595 110.280 58.765 112.540 ;
        RECT 59.135 111.970 67.175 112.140 ;
        RECT 67.345 110.910 67.515 111.910 ;
        RECT 59.135 110.680 67.175 110.850 ;
        RECT 67.855 110.280 68.025 112.540 ;
        RECT 58.595 110.110 68.025 110.280 ;
        RECT 74.480 111.960 74.650 114.220 ;
        RECT 75.020 113.650 83.060 113.820 ;
        RECT 83.230 112.590 83.400 113.590 ;
        RECT 75.020 112.360 83.060 112.530 ;
        RECT 83.740 111.960 83.910 114.220 ;
        RECT 84.585 113.260 84.755 115.520 ;
        RECT 85.125 114.950 93.165 115.120 ;
        RECT 93.380 113.890 93.550 114.890 ;
        RECT 85.125 113.660 93.165 113.830 ;
        RECT 93.895 113.260 94.065 115.520 ;
        RECT 84.585 113.090 94.065 113.260 ;
        RECT 74.480 111.790 83.910 111.960 ;
        RECT 48.480 109.360 57.910 109.530 ;
        RECT 48.480 107.100 48.650 109.360 ;
        RECT 49.020 108.790 57.060 108.960 ;
        RECT 57.230 107.730 57.400 108.730 ;
        RECT 49.020 107.500 57.060 107.670 ;
        RECT 57.740 107.100 57.910 109.360 ;
        RECT 48.480 106.930 57.910 107.100 ;
        RECT 48.480 104.670 48.650 106.930 ;
        RECT 49.020 106.360 57.060 106.530 ;
        RECT 57.230 105.300 57.400 106.300 ;
        RECT 49.020 105.070 57.060 105.240 ;
        RECT 57.740 104.670 57.910 106.930 ;
        RECT 48.480 104.500 57.910 104.670 ;
        RECT 58.580 109.550 68.060 109.720 ;
        RECT 58.580 107.320 58.750 109.550 ;
        RECT 59.120 108.980 67.160 109.150 ;
        RECT 67.375 107.920 67.545 108.920 ;
        RECT 59.120 107.690 67.160 107.860 ;
        RECT 67.890 107.320 68.060 109.550 ;
        RECT 58.580 107.120 68.060 107.320 ;
        RECT 58.580 104.920 58.750 107.120 ;
        RECT 59.120 106.580 67.160 106.750 ;
        RECT 67.375 105.520 67.545 106.520 ;
        RECT 59.120 105.290 67.160 105.460 ;
        RECT 67.890 104.920 68.060 107.120 ;
        RECT 58.580 104.720 68.060 104.920 ;
        RECT 48.480 104.450 57.810 104.500 ;
        RECT 35.180 104.110 40.660 104.280 ;
        RECT 17.030 103.060 19.630 103.065 ;
        RECT 6.200 102.890 11.230 103.060 ;
        RECT 6.200 93.750 6.370 102.890 ;
        RECT 7.000 102.375 8.000 102.545 ;
        RECT 6.770 94.120 6.940 102.160 ;
        RECT 8.060 94.120 8.230 102.160 ;
        RECT 8.630 93.750 8.800 102.890 ;
        RECT 9.430 102.375 10.430 102.545 ;
        RECT 9.200 94.120 9.370 102.160 ;
        RECT 10.490 94.120 10.660 102.160 ;
        RECT 11.060 93.750 11.230 102.890 ;
        RECT 6.200 93.580 11.230 93.750 ;
        RECT 11.600 102.840 14.200 103.010 ;
        RECT 11.600 93.750 11.770 102.840 ;
        RECT 12.400 102.330 13.400 102.500 ;
        RECT 12.170 94.120 12.340 102.160 ;
        RECT 13.460 94.120 13.630 102.160 ;
        RECT 14.030 93.750 14.200 102.840 ;
        RECT 11.600 93.580 14.200 93.750 ;
        RECT 14.600 102.895 19.630 103.060 ;
        RECT 14.600 102.890 17.200 102.895 ;
        RECT 14.600 93.750 14.770 102.890 ;
        RECT 15.400 102.375 16.400 102.545 ;
        RECT 15.170 94.120 15.340 102.160 ;
        RECT 16.460 94.120 16.630 102.160 ;
        RECT 17.030 93.755 17.200 102.890 ;
        RECT 17.830 102.380 18.830 102.550 ;
        RECT 17.600 94.125 17.770 102.165 ;
        RECT 18.890 94.125 19.060 102.165 ;
        RECT 19.460 93.755 19.630 102.895 ;
        RECT 17.030 93.750 19.630 93.755 ;
        RECT 14.600 93.585 19.630 93.750 ;
        RECT 20.010 102.855 22.610 103.025 ;
        RECT 20.010 93.765 20.180 102.855 ;
        RECT 20.810 102.345 21.810 102.515 ;
        RECT 20.580 94.135 20.750 102.175 ;
        RECT 21.870 94.135 22.040 102.175 ;
        RECT 22.440 93.765 22.610 102.855 ;
        RECT 20.010 93.595 22.610 93.765 ;
        RECT 23.000 102.890 32.795 103.060 ;
        RECT 23.000 93.750 23.170 102.890 ;
        RECT 23.800 102.375 24.800 102.545 ;
        RECT 23.570 94.120 23.740 102.160 ;
        RECT 24.860 94.120 25.030 102.160 ;
        RECT 25.400 93.750 25.600 102.890 ;
        RECT 26.200 102.375 27.200 102.545 ;
        RECT 25.970 94.120 26.140 102.160 ;
        RECT 27.260 94.120 27.430 102.160 ;
        RECT 27.800 93.750 28.000 102.890 ;
        RECT 28.600 102.375 29.600 102.545 ;
        RECT 28.370 94.120 28.540 102.160 ;
        RECT 29.660 94.120 29.830 102.160 ;
        RECT 30.195 93.750 30.400 102.890 ;
        RECT 30.995 102.375 31.995 102.545 ;
        RECT 30.765 94.120 30.935 102.160 ;
        RECT 32.055 94.120 32.225 102.160 ;
        RECT 32.625 98.480 32.795 102.890 ;
        RECT 35.180 102.350 35.350 104.110 ;
        RECT 35.720 103.540 39.760 103.710 ;
        RECT 39.975 102.980 40.145 103.480 ;
        RECT 35.720 102.750 39.760 102.920 ;
        RECT 40.490 102.350 40.660 104.110 ;
        RECT 35.180 102.180 40.660 102.350 ;
        RECT 33.200 100.560 42.800 100.730 ;
        RECT 33.200 99.050 33.370 100.560 ;
        RECT 34.000 100.050 42.000 100.220 ;
        RECT 33.770 99.420 33.940 99.880 ;
        RECT 42.060 99.420 42.230 99.880 ;
        RECT 42.630 99.050 42.800 100.560 ;
        RECT 33.200 98.880 42.800 99.050 ;
        RECT 32.625 98.310 42.300 98.480 ;
        RECT 32.625 96.750 32.870 98.310 ;
        RECT 33.500 97.795 41.500 97.965 ;
        RECT 33.270 97.120 33.440 97.580 ;
        RECT 41.560 97.120 41.730 97.580 ;
        RECT 42.130 96.750 42.300 98.310 ;
        RECT 32.625 96.580 42.300 96.750 ;
        RECT 32.625 93.750 32.795 96.580 ;
        RECT 14.600 93.580 17.200 93.585 ;
        RECT 23.000 93.580 32.795 93.750 ;
        RECT 33.200 96.010 42.630 96.180 ;
        RECT 33.200 93.750 33.370 96.010 ;
        RECT 33.740 95.440 41.780 95.610 ;
        RECT 41.950 94.380 42.120 95.380 ;
        RECT 33.740 94.150 41.780 94.320 ;
        RECT 42.460 93.750 42.630 96.010 ;
        RECT 48.480 95.190 48.650 104.450 ;
        RECT 49.020 103.880 50.060 104.050 ;
        RECT 50.230 95.820 50.400 103.820 ;
        RECT 49.020 95.590 50.060 95.760 ;
        RECT 50.740 95.190 50.950 104.450 ;
        RECT 51.320 103.880 52.360 104.050 ;
        RECT 52.530 95.820 52.700 103.820 ;
        RECT 51.320 95.590 52.360 95.760 ;
        RECT 53.040 95.190 53.250 104.450 ;
        RECT 53.620 103.880 54.660 104.050 ;
        RECT 54.830 95.820 55.000 103.820 ;
        RECT 53.620 95.590 54.660 95.760 ;
        RECT 55.340 95.190 55.550 104.450 ;
        RECT 55.920 103.880 56.960 104.050 ;
        RECT 48.480 95.020 55.550 95.190 ;
        RECT 33.200 93.580 42.630 93.750 ;
        RECT 6.180 92.810 28.220 92.910 ;
        RECT 6.180 92.740 42.800 92.810 ;
        RECT 6.180 83.650 6.350 92.740 ;
        RECT 6.980 92.230 7.980 92.400 ;
        RECT 6.750 84.020 6.920 92.060 ;
        RECT 8.040 84.020 8.210 92.060 ;
        RECT 8.610 83.650 8.780 92.740 ;
        RECT 9.410 92.230 10.410 92.400 ;
        RECT 9.180 84.020 9.350 92.060 ;
        RECT 10.470 84.020 10.640 92.060 ;
        RECT 11.040 83.650 11.210 92.740 ;
        RECT 11.840 92.230 12.840 92.400 ;
        RECT 11.610 84.020 11.780 92.060 ;
        RECT 12.900 84.020 13.070 92.060 ;
        RECT 13.470 83.650 13.640 92.740 ;
        RECT 14.270 92.230 15.270 92.400 ;
        RECT 14.040 84.020 14.210 92.060 ;
        RECT 15.330 84.020 15.500 92.060 ;
        RECT 15.900 83.650 16.070 92.740 ;
        RECT 16.700 92.230 17.700 92.400 ;
        RECT 16.470 84.020 16.640 92.060 ;
        RECT 17.760 84.020 17.930 92.060 ;
        RECT 18.330 83.650 18.500 92.740 ;
        RECT 19.130 92.230 20.130 92.400 ;
        RECT 18.900 84.020 19.070 92.060 ;
        RECT 20.190 84.020 20.360 92.060 ;
        RECT 20.760 83.650 20.930 92.740 ;
        RECT 21.560 92.230 22.560 92.400 ;
        RECT 21.330 84.020 21.500 92.060 ;
        RECT 22.620 84.020 22.790 92.060 ;
        RECT 23.190 83.650 23.360 92.740 ;
        RECT 23.990 92.230 24.990 92.400 ;
        RECT 23.760 84.020 23.930 92.060 ;
        RECT 25.050 84.020 25.220 92.060 ;
        RECT 25.620 83.650 25.790 92.740 ;
        RECT 28.050 92.640 42.800 92.740 ;
        RECT 26.420 92.230 27.420 92.400 ;
        RECT 26.190 84.020 26.360 92.060 ;
        RECT 27.480 84.020 27.650 92.060 ;
        RECT 28.050 90.550 28.270 92.640 ;
        RECT 28.900 92.130 42.000 92.300 ;
        RECT 28.670 90.920 28.840 91.960 ;
        RECT 42.060 90.920 42.230 91.960 ;
        RECT 42.630 90.550 42.800 92.640 ;
        RECT 28.050 90.380 42.800 90.550 ;
        RECT 28.050 90.340 37.700 90.380 ;
        RECT 28.050 88.250 28.270 90.340 ;
        RECT 28.900 89.830 36.900 90.000 ;
        RECT 28.670 88.620 28.840 89.660 ;
        RECT 36.960 88.620 37.130 89.660 ;
        RECT 37.530 88.250 37.700 90.340 ;
        RECT 55.380 90.090 55.550 95.020 ;
        RECT 57.130 90.720 57.300 103.820 ;
        RECT 55.920 90.490 56.960 90.660 ;
        RECT 57.640 90.090 57.810 104.450 ;
        RECT 58.580 102.525 58.750 104.720 ;
        RECT 59.120 104.180 67.160 104.350 ;
        RECT 67.375 103.120 67.545 104.120 ;
        RECT 59.120 102.890 67.160 103.060 ;
        RECT 67.890 102.525 68.060 104.720 ;
        RECT 58.580 102.320 68.060 102.525 ;
        RECT 58.580 100.095 58.750 102.320 ;
        RECT 59.120 101.785 67.160 101.955 ;
        RECT 67.375 100.725 67.545 101.725 ;
        RECT 59.120 100.495 67.160 100.665 ;
        RECT 67.890 100.095 68.060 102.320 ;
        RECT 58.580 99.925 68.060 100.095 ;
        RECT 74.480 109.530 74.650 111.790 ;
        RECT 75.020 111.220 83.060 111.390 ;
        RECT 83.230 110.160 83.400 111.160 ;
        RECT 75.020 109.930 83.060 110.100 ;
        RECT 83.740 109.530 83.910 111.790 ;
        RECT 84.595 112.540 94.025 112.710 ;
        RECT 84.595 110.280 84.765 112.540 ;
        RECT 85.135 111.970 93.175 112.140 ;
        RECT 93.345 110.910 93.515 111.910 ;
        RECT 85.135 110.680 93.175 110.850 ;
        RECT 93.855 110.280 94.025 112.540 ;
        RECT 84.595 110.110 94.025 110.280 ;
        RECT 74.480 109.360 83.910 109.530 ;
        RECT 74.480 107.100 74.650 109.360 ;
        RECT 75.020 108.790 83.060 108.960 ;
        RECT 83.230 107.730 83.400 108.730 ;
        RECT 75.020 107.500 83.060 107.670 ;
        RECT 83.740 107.100 83.910 109.360 ;
        RECT 74.480 106.930 83.910 107.100 ;
        RECT 74.480 104.670 74.650 106.930 ;
        RECT 75.020 106.360 83.060 106.530 ;
        RECT 83.230 105.300 83.400 106.300 ;
        RECT 75.020 105.070 83.060 105.240 ;
        RECT 83.740 104.670 83.910 106.930 ;
        RECT 74.480 104.500 83.910 104.670 ;
        RECT 84.580 109.550 94.060 109.720 ;
        RECT 84.580 107.320 84.750 109.550 ;
        RECT 85.120 108.980 93.160 109.150 ;
        RECT 93.375 107.920 93.545 108.920 ;
        RECT 85.120 107.690 93.160 107.860 ;
        RECT 93.890 107.320 94.060 109.550 ;
        RECT 84.580 107.120 94.060 107.320 ;
        RECT 84.580 104.920 84.750 107.120 ;
        RECT 85.120 106.580 93.160 106.750 ;
        RECT 93.375 105.520 93.545 106.520 ;
        RECT 85.120 105.290 93.160 105.460 ;
        RECT 93.890 104.920 94.060 107.120 ;
        RECT 84.580 104.720 94.060 104.920 ;
        RECT 74.480 104.450 83.810 104.500 ;
        RECT 61.580 99.850 63.480 99.925 ;
        RECT 58.580 99.350 61.180 99.520 ;
        RECT 58.580 90.260 58.750 99.350 ;
        RECT 59.150 90.940 59.320 98.980 ;
        RECT 60.440 90.940 60.610 98.980 ;
        RECT 59.380 90.600 60.380 90.770 ;
        RECT 61.010 90.260 61.180 99.350 ;
        RECT 61.580 90.590 61.750 99.850 ;
        RECT 62.120 99.280 62.580 99.450 ;
        RECT 62.795 91.220 62.965 99.220 ;
        RECT 62.120 90.990 62.580 91.160 ;
        RECT 63.310 90.590 63.480 99.850 ;
        RECT 61.580 90.420 63.480 90.590 ;
        RECT 63.880 99.350 65.730 99.520 ;
        RECT 58.580 90.090 61.180 90.260 ;
        RECT 63.880 90.090 64.050 99.350 ;
        RECT 64.420 98.780 64.880 98.950 ;
        RECT 65.050 90.720 65.220 98.720 ;
        RECT 64.420 90.490 64.880 90.660 ;
        RECT 65.560 90.090 65.730 99.350 ;
        RECT 67.180 97.490 69.280 97.660 ;
        RECT 67.180 92.350 67.350 97.490 ;
        RECT 67.750 93.080 67.920 97.120 ;
        RECT 68.540 93.080 68.710 97.120 ;
        RECT 67.980 92.695 68.480 92.865 ;
        RECT 69.110 92.350 69.280 97.490 ;
        RECT 74.480 95.190 74.650 104.450 ;
        RECT 75.020 103.880 76.060 104.050 ;
        RECT 76.230 95.820 76.400 103.820 ;
        RECT 75.020 95.590 76.060 95.760 ;
        RECT 76.740 95.190 76.950 104.450 ;
        RECT 77.320 103.880 78.360 104.050 ;
        RECT 78.530 95.820 78.700 103.820 ;
        RECT 77.320 95.590 78.360 95.760 ;
        RECT 79.040 95.190 79.250 104.450 ;
        RECT 79.620 103.880 80.660 104.050 ;
        RECT 80.830 95.820 81.000 103.820 ;
        RECT 79.620 95.590 80.660 95.760 ;
        RECT 81.340 95.190 81.550 104.450 ;
        RECT 81.920 103.880 82.960 104.050 ;
        RECT 74.480 95.020 81.550 95.190 ;
        RECT 67.180 92.180 69.280 92.350 ;
        RECT 55.380 89.920 57.810 90.090 ;
        RECT 63.880 89.920 65.730 90.090 ;
        RECT 81.380 90.090 81.550 95.020 ;
        RECT 83.130 90.720 83.300 103.820 ;
        RECT 81.920 90.490 82.960 90.660 ;
        RECT 83.640 90.090 83.810 104.450 ;
        RECT 84.580 102.525 84.750 104.720 ;
        RECT 85.120 104.180 93.160 104.350 ;
        RECT 93.375 103.120 93.545 104.120 ;
        RECT 85.120 102.890 93.160 103.060 ;
        RECT 93.890 102.525 94.060 104.720 ;
        RECT 84.580 102.320 94.060 102.525 ;
        RECT 84.580 100.095 84.750 102.320 ;
        RECT 85.120 101.785 93.160 101.955 ;
        RECT 93.375 100.725 93.545 101.725 ;
        RECT 85.120 100.495 93.160 100.665 ;
        RECT 93.890 100.095 94.060 102.320 ;
        RECT 84.580 99.925 94.060 100.095 ;
        RECT 87.580 99.850 89.480 99.925 ;
        RECT 84.580 99.350 87.180 99.520 ;
        RECT 84.580 90.260 84.750 99.350 ;
        RECT 85.150 90.940 85.320 98.980 ;
        RECT 86.440 90.940 86.610 98.980 ;
        RECT 85.380 90.600 86.380 90.770 ;
        RECT 87.010 90.260 87.180 99.350 ;
        RECT 87.580 90.590 87.750 99.850 ;
        RECT 88.120 99.280 88.580 99.450 ;
        RECT 88.795 91.220 88.965 99.220 ;
        RECT 88.120 90.990 88.580 91.160 ;
        RECT 89.310 90.590 89.480 99.850 ;
        RECT 87.580 90.420 89.480 90.590 ;
        RECT 89.880 99.350 91.730 99.520 ;
        RECT 84.580 90.090 87.180 90.260 ;
        RECT 89.880 90.090 90.050 99.350 ;
        RECT 90.420 98.780 90.880 98.950 ;
        RECT 91.050 90.720 91.220 98.720 ;
        RECT 90.420 90.490 90.880 90.660 ;
        RECT 91.560 90.090 91.730 99.350 ;
        RECT 93.180 97.490 95.280 97.660 ;
        RECT 93.180 92.350 93.350 97.490 ;
        RECT 93.750 93.080 93.920 97.120 ;
        RECT 94.540 93.080 94.710 97.120 ;
        RECT 93.980 92.695 94.480 92.865 ;
        RECT 95.110 92.350 95.280 97.490 ;
        RECT 93.180 92.180 95.280 92.350 ;
        RECT 81.380 89.920 83.810 90.090 ;
        RECT 89.880 89.920 91.730 90.090 ;
        RECT 28.050 88.040 37.700 88.250 ;
        RECT 28.050 85.950 28.270 88.040 ;
        RECT 28.900 87.530 36.900 87.700 ;
        RECT 28.670 86.320 28.840 87.360 ;
        RECT 36.960 86.320 37.130 87.360 ;
        RECT 37.530 85.950 37.700 88.040 ;
        RECT 28.050 85.740 37.700 85.950 ;
        RECT 28.050 83.650 28.270 85.740 ;
        RECT 28.900 85.230 36.900 85.400 ;
        RECT 28.670 84.020 28.840 85.060 ;
        RECT 36.960 84.020 37.130 85.060 ;
        RECT 37.530 83.650 37.700 85.740 ;
        RECT 6.180 83.480 37.700 83.650 ;
        RECT 48.480 84.370 57.910 84.540 ;
        RECT 48.480 82.110 48.650 84.370 ;
        RECT 49.020 83.800 57.060 83.970 ;
        RECT 57.230 82.740 57.400 83.740 ;
        RECT 49.020 82.510 57.060 82.680 ;
        RECT 57.740 82.110 57.910 84.370 ;
        RECT 48.480 81.940 57.910 82.110 ;
        RECT 48.480 79.680 48.650 81.940 ;
        RECT 49.020 81.370 57.060 81.540 ;
        RECT 57.230 80.310 57.400 81.310 ;
        RECT 49.020 80.080 57.060 80.250 ;
        RECT 57.740 79.680 57.910 81.940 ;
        RECT 48.480 79.510 57.910 79.680 ;
        RECT 35.180 78.110 40.660 78.280 ;
        RECT 17.030 77.060 19.630 77.065 ;
        RECT 6.200 76.890 11.230 77.060 ;
        RECT 6.200 67.750 6.370 76.890 ;
        RECT 7.000 76.375 8.000 76.545 ;
        RECT 6.770 68.120 6.940 76.160 ;
        RECT 8.060 68.120 8.230 76.160 ;
        RECT 8.630 67.750 8.800 76.890 ;
        RECT 9.430 76.375 10.430 76.545 ;
        RECT 9.200 68.120 9.370 76.160 ;
        RECT 10.490 68.120 10.660 76.160 ;
        RECT 11.060 67.750 11.230 76.890 ;
        RECT 6.200 67.580 11.230 67.750 ;
        RECT 11.600 76.840 14.200 77.010 ;
        RECT 11.600 67.750 11.770 76.840 ;
        RECT 12.400 76.330 13.400 76.500 ;
        RECT 12.170 68.120 12.340 76.160 ;
        RECT 13.460 68.120 13.630 76.160 ;
        RECT 14.030 67.750 14.200 76.840 ;
        RECT 11.600 67.580 14.200 67.750 ;
        RECT 14.600 76.895 19.630 77.060 ;
        RECT 14.600 76.890 17.200 76.895 ;
        RECT 14.600 67.750 14.770 76.890 ;
        RECT 15.400 76.375 16.400 76.545 ;
        RECT 15.170 68.120 15.340 76.160 ;
        RECT 16.460 68.120 16.630 76.160 ;
        RECT 17.030 67.755 17.200 76.890 ;
        RECT 17.830 76.380 18.830 76.550 ;
        RECT 17.600 68.125 17.770 76.165 ;
        RECT 18.890 68.125 19.060 76.165 ;
        RECT 19.460 67.755 19.630 76.895 ;
        RECT 17.030 67.750 19.630 67.755 ;
        RECT 14.600 67.585 19.630 67.750 ;
        RECT 20.010 76.855 22.610 77.025 ;
        RECT 20.010 67.765 20.180 76.855 ;
        RECT 20.810 76.345 21.810 76.515 ;
        RECT 20.580 68.135 20.750 76.175 ;
        RECT 21.870 68.135 22.040 76.175 ;
        RECT 22.440 67.765 22.610 76.855 ;
        RECT 20.010 67.595 22.610 67.765 ;
        RECT 23.000 76.890 32.795 77.060 ;
        RECT 23.000 67.750 23.170 76.890 ;
        RECT 23.800 76.375 24.800 76.545 ;
        RECT 23.570 68.120 23.740 76.160 ;
        RECT 24.860 68.120 25.030 76.160 ;
        RECT 25.400 67.750 25.600 76.890 ;
        RECT 26.200 76.375 27.200 76.545 ;
        RECT 25.970 68.120 26.140 76.160 ;
        RECT 27.260 68.120 27.430 76.160 ;
        RECT 27.800 67.750 28.000 76.890 ;
        RECT 28.600 76.375 29.600 76.545 ;
        RECT 28.370 68.120 28.540 76.160 ;
        RECT 29.660 68.120 29.830 76.160 ;
        RECT 30.195 67.750 30.400 76.890 ;
        RECT 30.995 76.375 31.995 76.545 ;
        RECT 30.765 68.120 30.935 76.160 ;
        RECT 32.055 68.120 32.225 76.160 ;
        RECT 32.625 72.480 32.795 76.890 ;
        RECT 35.180 76.350 35.350 78.110 ;
        RECT 35.720 77.540 39.760 77.710 ;
        RECT 39.975 76.980 40.145 77.480 ;
        RECT 35.720 76.750 39.760 76.920 ;
        RECT 40.490 76.350 40.660 78.110 ;
        RECT 35.180 76.180 40.660 76.350 ;
        RECT 48.480 77.250 48.650 79.510 ;
        RECT 49.020 78.940 57.060 79.110 ;
        RECT 57.230 77.880 57.400 78.880 ;
        RECT 49.020 77.650 57.060 77.820 ;
        RECT 57.740 77.250 57.910 79.510 ;
        RECT 58.580 84.350 68.060 84.520 ;
        RECT 58.580 82.090 58.750 84.350 ;
        RECT 59.120 83.780 67.160 83.950 ;
        RECT 67.375 82.720 67.545 83.720 ;
        RECT 59.120 82.490 67.160 82.660 ;
        RECT 67.890 82.090 68.060 84.350 ;
        RECT 58.580 81.920 68.060 82.090 ;
        RECT 58.580 79.660 58.750 81.920 ;
        RECT 59.120 81.350 67.160 81.520 ;
        RECT 67.375 80.290 67.545 81.290 ;
        RECT 59.120 80.060 67.160 80.230 ;
        RECT 67.890 79.660 68.060 81.920 ;
        RECT 58.580 79.490 68.060 79.660 ;
        RECT 74.480 84.370 83.910 84.540 ;
        RECT 74.480 82.110 74.650 84.370 ;
        RECT 75.020 83.800 83.060 83.970 ;
        RECT 83.230 82.740 83.400 83.740 ;
        RECT 75.020 82.510 83.060 82.680 ;
        RECT 83.740 82.110 83.910 84.370 ;
        RECT 74.480 81.940 83.910 82.110 ;
        RECT 74.480 79.680 74.650 81.940 ;
        RECT 75.020 81.370 83.060 81.540 ;
        RECT 83.230 80.310 83.400 81.310 ;
        RECT 75.020 80.080 83.060 80.250 ;
        RECT 83.740 79.680 83.910 81.940 ;
        RECT 74.480 79.510 83.910 79.680 ;
        RECT 48.480 77.080 57.910 77.250 ;
        RECT 48.480 74.820 48.650 77.080 ;
        RECT 49.020 76.510 57.060 76.680 ;
        RECT 57.230 75.450 57.400 76.450 ;
        RECT 49.020 75.220 57.060 75.390 ;
        RECT 57.740 74.820 57.910 77.080 ;
        RECT 58.580 78.950 68.010 79.120 ;
        RECT 58.580 76.690 58.750 78.950 ;
        RECT 59.120 78.380 67.160 78.550 ;
        RECT 67.330 77.320 67.500 78.320 ;
        RECT 59.120 77.090 67.160 77.260 ;
        RECT 67.840 76.690 68.010 78.950 ;
        RECT 58.580 76.520 68.010 76.690 ;
        RECT 74.480 77.250 74.650 79.510 ;
        RECT 75.020 78.940 83.060 79.110 ;
        RECT 83.230 77.880 83.400 78.880 ;
        RECT 75.020 77.650 83.060 77.820 ;
        RECT 83.740 77.250 83.910 79.510 ;
        RECT 84.580 84.350 94.060 84.520 ;
        RECT 84.580 82.090 84.750 84.350 ;
        RECT 85.120 83.780 93.160 83.950 ;
        RECT 93.375 82.720 93.545 83.720 ;
        RECT 85.120 82.490 93.160 82.660 ;
        RECT 93.890 82.090 94.060 84.350 ;
        RECT 84.580 81.920 94.060 82.090 ;
        RECT 84.580 79.660 84.750 81.920 ;
        RECT 85.120 81.350 93.160 81.520 ;
        RECT 93.375 80.290 93.545 81.290 ;
        RECT 85.120 80.060 93.160 80.230 ;
        RECT 93.890 79.660 94.060 81.920 ;
        RECT 84.580 79.490 94.060 79.660 ;
        RECT 74.480 77.080 83.910 77.250 ;
        RECT 33.200 74.560 42.800 74.730 ;
        RECT 33.200 73.050 33.370 74.560 ;
        RECT 34.000 74.050 42.000 74.220 ;
        RECT 33.770 73.420 33.940 73.880 ;
        RECT 42.060 73.420 42.230 73.880 ;
        RECT 42.630 73.050 42.800 74.560 ;
        RECT 33.200 72.880 42.800 73.050 ;
        RECT 48.480 74.650 57.910 74.820 ;
        RECT 32.625 72.310 42.300 72.480 ;
        RECT 32.625 70.750 32.870 72.310 ;
        RECT 33.500 71.795 41.500 71.965 ;
        RECT 33.270 71.120 33.440 71.580 ;
        RECT 41.560 71.120 41.730 71.580 ;
        RECT 42.130 70.750 42.300 72.310 ;
        RECT 32.625 70.580 42.300 70.750 ;
        RECT 48.480 72.390 48.650 74.650 ;
        RECT 49.020 74.080 57.060 74.250 ;
        RECT 57.230 73.020 57.400 74.020 ;
        RECT 49.020 72.790 57.060 72.960 ;
        RECT 57.740 72.390 57.910 74.650 ;
        RECT 58.580 75.950 68.060 76.120 ;
        RECT 58.580 73.690 58.750 75.950 ;
        RECT 59.120 75.380 67.160 75.550 ;
        RECT 67.375 74.320 67.545 75.320 ;
        RECT 59.120 74.090 67.160 74.260 ;
        RECT 67.890 73.690 68.060 75.950 ;
        RECT 74.480 74.820 74.650 77.080 ;
        RECT 75.020 76.510 83.060 76.680 ;
        RECT 83.230 75.450 83.400 76.450 ;
        RECT 75.020 75.220 83.060 75.390 ;
        RECT 83.740 74.820 83.910 77.080 ;
        RECT 84.580 78.950 94.010 79.120 ;
        RECT 84.580 76.690 84.750 78.950 ;
        RECT 85.120 78.380 93.160 78.550 ;
        RECT 93.330 77.320 93.500 78.320 ;
        RECT 85.120 77.090 93.160 77.260 ;
        RECT 93.840 76.690 94.010 78.950 ;
        RECT 84.580 76.520 94.010 76.690 ;
        RECT 74.480 74.650 83.910 74.820 ;
        RECT 58.580 73.520 68.065 73.690 ;
        RECT 48.480 72.220 57.910 72.390 ;
        RECT 32.625 67.750 32.795 70.580 ;
        RECT 14.600 67.580 17.200 67.585 ;
        RECT 23.000 67.580 32.795 67.750 ;
        RECT 33.200 70.010 42.630 70.180 ;
        RECT 33.200 67.750 33.370 70.010 ;
        RECT 33.740 69.440 41.780 69.610 ;
        RECT 41.950 68.380 42.120 69.380 ;
        RECT 33.740 68.150 41.780 68.320 ;
        RECT 42.460 67.750 42.630 70.010 ;
        RECT 33.200 67.580 42.630 67.750 ;
        RECT 48.480 69.960 48.650 72.220 ;
        RECT 49.020 71.650 57.060 71.820 ;
        RECT 57.230 70.590 57.400 71.590 ;
        RECT 49.020 70.360 57.060 70.530 ;
        RECT 57.740 69.960 57.910 72.220 ;
        RECT 58.585 71.260 58.755 73.520 ;
        RECT 59.125 72.950 67.165 73.120 ;
        RECT 67.380 71.890 67.550 72.890 ;
        RECT 59.125 71.660 67.165 71.830 ;
        RECT 67.895 71.260 68.065 73.520 ;
        RECT 58.585 71.090 68.065 71.260 ;
        RECT 74.480 72.390 74.650 74.650 ;
        RECT 75.020 74.080 83.060 74.250 ;
        RECT 83.230 73.020 83.400 74.020 ;
        RECT 75.020 72.790 83.060 72.960 ;
        RECT 83.740 72.390 83.910 74.650 ;
        RECT 84.580 75.950 94.060 76.120 ;
        RECT 84.580 73.690 84.750 75.950 ;
        RECT 85.120 75.380 93.160 75.550 ;
        RECT 93.375 74.320 93.545 75.320 ;
        RECT 85.120 74.090 93.160 74.260 ;
        RECT 93.890 73.690 94.060 75.950 ;
        RECT 84.580 73.520 94.065 73.690 ;
        RECT 74.480 72.220 83.910 72.390 ;
        RECT 48.480 69.790 57.910 69.960 ;
        RECT 48.480 67.530 48.650 69.790 ;
        RECT 49.020 69.220 57.060 69.390 ;
        RECT 57.230 68.160 57.400 69.160 ;
        RECT 49.020 67.930 57.060 68.100 ;
        RECT 57.740 67.530 57.910 69.790 ;
        RECT 58.595 70.540 68.025 70.710 ;
        RECT 58.595 68.280 58.765 70.540 ;
        RECT 59.135 69.970 67.175 70.140 ;
        RECT 67.345 68.910 67.515 69.910 ;
        RECT 59.135 68.680 67.175 68.850 ;
        RECT 67.855 68.280 68.025 70.540 ;
        RECT 58.595 68.110 68.025 68.280 ;
        RECT 74.480 69.960 74.650 72.220 ;
        RECT 75.020 71.650 83.060 71.820 ;
        RECT 83.230 70.590 83.400 71.590 ;
        RECT 75.020 70.360 83.060 70.530 ;
        RECT 83.740 69.960 83.910 72.220 ;
        RECT 84.585 71.260 84.755 73.520 ;
        RECT 85.125 72.950 93.165 73.120 ;
        RECT 93.380 71.890 93.550 72.890 ;
        RECT 85.125 71.660 93.165 71.830 ;
        RECT 93.895 71.260 94.065 73.520 ;
        RECT 84.585 71.090 94.065 71.260 ;
        RECT 74.480 69.790 83.910 69.960 ;
        RECT 48.480 67.360 57.910 67.530 ;
        RECT 6.180 66.810 28.220 66.910 ;
        RECT 6.180 66.740 42.800 66.810 ;
        RECT 6.180 57.650 6.350 66.740 ;
        RECT 6.980 66.230 7.980 66.400 ;
        RECT 6.750 58.020 6.920 66.060 ;
        RECT 8.040 58.020 8.210 66.060 ;
        RECT 8.610 57.650 8.780 66.740 ;
        RECT 9.410 66.230 10.410 66.400 ;
        RECT 9.180 58.020 9.350 66.060 ;
        RECT 10.470 58.020 10.640 66.060 ;
        RECT 11.040 57.650 11.210 66.740 ;
        RECT 11.840 66.230 12.840 66.400 ;
        RECT 11.610 58.020 11.780 66.060 ;
        RECT 12.900 58.020 13.070 66.060 ;
        RECT 13.470 57.650 13.640 66.740 ;
        RECT 14.270 66.230 15.270 66.400 ;
        RECT 14.040 58.020 14.210 66.060 ;
        RECT 15.330 58.020 15.500 66.060 ;
        RECT 15.900 57.650 16.070 66.740 ;
        RECT 16.700 66.230 17.700 66.400 ;
        RECT 16.470 58.020 16.640 66.060 ;
        RECT 17.760 58.020 17.930 66.060 ;
        RECT 18.330 57.650 18.500 66.740 ;
        RECT 19.130 66.230 20.130 66.400 ;
        RECT 18.900 58.020 19.070 66.060 ;
        RECT 20.190 58.020 20.360 66.060 ;
        RECT 20.760 57.650 20.930 66.740 ;
        RECT 21.560 66.230 22.560 66.400 ;
        RECT 21.330 58.020 21.500 66.060 ;
        RECT 22.620 58.020 22.790 66.060 ;
        RECT 23.190 57.650 23.360 66.740 ;
        RECT 23.990 66.230 24.990 66.400 ;
        RECT 23.760 58.020 23.930 66.060 ;
        RECT 25.050 58.020 25.220 66.060 ;
        RECT 25.620 57.650 25.790 66.740 ;
        RECT 28.050 66.640 42.800 66.740 ;
        RECT 26.420 66.230 27.420 66.400 ;
        RECT 26.190 58.020 26.360 66.060 ;
        RECT 27.480 58.020 27.650 66.060 ;
        RECT 28.050 64.550 28.270 66.640 ;
        RECT 28.900 66.130 42.000 66.300 ;
        RECT 28.670 64.920 28.840 65.960 ;
        RECT 42.060 64.920 42.230 65.960 ;
        RECT 42.630 64.550 42.800 66.640 ;
        RECT 28.050 64.380 42.800 64.550 ;
        RECT 48.480 65.100 48.650 67.360 ;
        RECT 49.020 66.790 57.060 66.960 ;
        RECT 57.230 65.730 57.400 66.730 ;
        RECT 49.020 65.500 57.060 65.670 ;
        RECT 57.740 65.100 57.910 67.360 ;
        RECT 48.480 64.930 57.910 65.100 ;
        RECT 28.050 64.340 37.700 64.380 ;
        RECT 28.050 62.250 28.270 64.340 ;
        RECT 28.900 63.830 36.900 64.000 ;
        RECT 28.670 62.620 28.840 63.660 ;
        RECT 36.960 62.620 37.130 63.660 ;
        RECT 37.530 62.250 37.700 64.340 ;
        RECT 28.050 62.040 37.700 62.250 ;
        RECT 28.050 59.950 28.270 62.040 ;
        RECT 28.900 61.530 36.900 61.700 ;
        RECT 28.670 60.320 28.840 61.360 ;
        RECT 36.960 60.320 37.130 61.360 ;
        RECT 37.530 59.950 37.700 62.040 ;
        RECT 28.050 59.740 37.700 59.950 ;
        RECT 28.050 57.650 28.270 59.740 ;
        RECT 28.900 59.230 36.900 59.400 ;
        RECT 28.670 58.020 28.840 59.060 ;
        RECT 36.960 58.020 37.130 59.060 ;
        RECT 37.530 57.650 37.700 59.740 ;
        RECT 6.180 57.480 37.700 57.650 ;
        RECT 48.480 62.670 48.650 64.930 ;
        RECT 49.020 64.360 57.060 64.530 ;
        RECT 57.230 63.300 57.400 64.300 ;
        RECT 49.020 63.070 57.060 63.240 ;
        RECT 57.740 62.670 57.910 64.930 ;
        RECT 48.480 62.500 57.910 62.670 ;
        RECT 58.580 67.550 68.060 67.720 ;
        RECT 58.580 65.320 58.750 67.550 ;
        RECT 59.120 66.980 67.160 67.150 ;
        RECT 67.375 65.920 67.545 66.920 ;
        RECT 59.120 65.690 67.160 65.860 ;
        RECT 67.890 65.320 68.060 67.550 ;
        RECT 58.580 65.120 68.060 65.320 ;
        RECT 58.580 62.920 58.750 65.120 ;
        RECT 59.120 64.580 67.160 64.750 ;
        RECT 67.375 63.520 67.545 64.520 ;
        RECT 59.120 63.290 67.160 63.460 ;
        RECT 67.890 62.920 68.060 65.120 ;
        RECT 58.580 62.720 68.060 62.920 ;
        RECT 48.480 62.450 57.810 62.500 ;
        RECT 48.480 53.190 48.650 62.450 ;
        RECT 49.020 61.880 50.060 62.050 ;
        RECT 50.230 53.820 50.400 61.820 ;
        RECT 49.020 53.590 50.060 53.760 ;
        RECT 50.740 53.190 50.950 62.450 ;
        RECT 51.320 61.880 52.360 62.050 ;
        RECT 52.530 53.820 52.700 61.820 ;
        RECT 51.320 53.590 52.360 53.760 ;
        RECT 53.040 53.190 53.250 62.450 ;
        RECT 53.620 61.880 54.660 62.050 ;
        RECT 54.830 53.820 55.000 61.820 ;
        RECT 53.620 53.590 54.660 53.760 ;
        RECT 55.340 53.190 55.550 62.450 ;
        RECT 55.920 61.880 56.960 62.050 ;
        RECT 48.480 53.020 55.550 53.190 ;
        RECT 35.180 52.110 40.660 52.280 ;
        RECT 17.030 51.060 19.630 51.065 ;
        RECT 6.200 50.890 11.230 51.060 ;
        RECT 6.200 41.750 6.370 50.890 ;
        RECT 7.000 50.375 8.000 50.545 ;
        RECT 6.770 42.120 6.940 50.160 ;
        RECT 8.060 42.120 8.230 50.160 ;
        RECT 8.630 41.750 8.800 50.890 ;
        RECT 9.430 50.375 10.430 50.545 ;
        RECT 9.200 42.120 9.370 50.160 ;
        RECT 10.490 42.120 10.660 50.160 ;
        RECT 11.060 41.750 11.230 50.890 ;
        RECT 6.200 41.580 11.230 41.750 ;
        RECT 11.600 50.840 14.200 51.010 ;
        RECT 11.600 41.750 11.770 50.840 ;
        RECT 12.400 50.330 13.400 50.500 ;
        RECT 12.170 42.120 12.340 50.160 ;
        RECT 13.460 42.120 13.630 50.160 ;
        RECT 14.030 41.750 14.200 50.840 ;
        RECT 11.600 41.580 14.200 41.750 ;
        RECT 14.600 50.895 19.630 51.060 ;
        RECT 14.600 50.890 17.200 50.895 ;
        RECT 14.600 41.750 14.770 50.890 ;
        RECT 15.400 50.375 16.400 50.545 ;
        RECT 15.170 42.120 15.340 50.160 ;
        RECT 16.460 42.120 16.630 50.160 ;
        RECT 17.030 41.755 17.200 50.890 ;
        RECT 17.830 50.380 18.830 50.550 ;
        RECT 17.600 42.125 17.770 50.165 ;
        RECT 18.890 42.125 19.060 50.165 ;
        RECT 19.460 41.755 19.630 50.895 ;
        RECT 17.030 41.750 19.630 41.755 ;
        RECT 14.600 41.585 19.630 41.750 ;
        RECT 20.010 50.855 22.610 51.025 ;
        RECT 20.010 41.765 20.180 50.855 ;
        RECT 20.810 50.345 21.810 50.515 ;
        RECT 20.580 42.135 20.750 50.175 ;
        RECT 21.870 42.135 22.040 50.175 ;
        RECT 22.440 41.765 22.610 50.855 ;
        RECT 20.010 41.595 22.610 41.765 ;
        RECT 23.000 50.890 32.795 51.060 ;
        RECT 23.000 41.750 23.170 50.890 ;
        RECT 23.800 50.375 24.800 50.545 ;
        RECT 23.570 42.120 23.740 50.160 ;
        RECT 24.860 42.120 25.030 50.160 ;
        RECT 25.400 41.750 25.600 50.890 ;
        RECT 26.200 50.375 27.200 50.545 ;
        RECT 25.970 42.120 26.140 50.160 ;
        RECT 27.260 42.120 27.430 50.160 ;
        RECT 27.800 41.750 28.000 50.890 ;
        RECT 28.600 50.375 29.600 50.545 ;
        RECT 28.370 42.120 28.540 50.160 ;
        RECT 29.660 42.120 29.830 50.160 ;
        RECT 30.195 41.750 30.400 50.890 ;
        RECT 30.995 50.375 31.995 50.545 ;
        RECT 30.765 42.120 30.935 50.160 ;
        RECT 32.055 42.120 32.225 50.160 ;
        RECT 32.625 46.480 32.795 50.890 ;
        RECT 35.180 50.350 35.350 52.110 ;
        RECT 35.720 51.540 39.760 51.710 ;
        RECT 39.975 50.980 40.145 51.480 ;
        RECT 35.720 50.750 39.760 50.920 ;
        RECT 40.490 50.350 40.660 52.110 ;
        RECT 35.180 50.180 40.660 50.350 ;
        RECT 33.200 48.560 42.800 48.730 ;
        RECT 33.200 47.050 33.370 48.560 ;
        RECT 34.000 48.050 42.000 48.220 ;
        RECT 33.770 47.420 33.940 47.880 ;
        RECT 42.060 47.420 42.230 47.880 ;
        RECT 42.630 47.050 42.800 48.560 ;
        RECT 55.380 48.090 55.550 53.020 ;
        RECT 57.130 48.720 57.300 61.820 ;
        RECT 55.920 48.490 56.960 48.660 ;
        RECT 57.640 48.090 57.810 62.450 ;
        RECT 58.580 60.525 58.750 62.720 ;
        RECT 59.120 62.180 67.160 62.350 ;
        RECT 67.375 61.120 67.545 62.120 ;
        RECT 59.120 60.890 67.160 61.060 ;
        RECT 67.890 60.525 68.060 62.720 ;
        RECT 58.580 60.320 68.060 60.525 ;
        RECT 58.580 58.095 58.750 60.320 ;
        RECT 59.120 59.785 67.160 59.955 ;
        RECT 67.375 58.725 67.545 59.725 ;
        RECT 59.120 58.495 67.160 58.665 ;
        RECT 67.890 58.095 68.060 60.320 ;
        RECT 58.580 57.925 68.060 58.095 ;
        RECT 74.480 67.530 74.650 69.790 ;
        RECT 75.020 69.220 83.060 69.390 ;
        RECT 83.230 68.160 83.400 69.160 ;
        RECT 75.020 67.930 83.060 68.100 ;
        RECT 83.740 67.530 83.910 69.790 ;
        RECT 84.595 70.540 94.025 70.710 ;
        RECT 84.595 68.280 84.765 70.540 ;
        RECT 85.135 69.970 93.175 70.140 ;
        RECT 93.345 68.910 93.515 69.910 ;
        RECT 85.135 68.680 93.175 68.850 ;
        RECT 93.855 68.280 94.025 70.540 ;
        RECT 84.595 68.110 94.025 68.280 ;
        RECT 74.480 67.360 83.910 67.530 ;
        RECT 74.480 65.100 74.650 67.360 ;
        RECT 75.020 66.790 83.060 66.960 ;
        RECT 83.230 65.730 83.400 66.730 ;
        RECT 75.020 65.500 83.060 65.670 ;
        RECT 83.740 65.100 83.910 67.360 ;
        RECT 74.480 64.930 83.910 65.100 ;
        RECT 74.480 62.670 74.650 64.930 ;
        RECT 75.020 64.360 83.060 64.530 ;
        RECT 83.230 63.300 83.400 64.300 ;
        RECT 75.020 63.070 83.060 63.240 ;
        RECT 83.740 62.670 83.910 64.930 ;
        RECT 74.480 62.500 83.910 62.670 ;
        RECT 84.580 67.550 94.060 67.720 ;
        RECT 84.580 65.320 84.750 67.550 ;
        RECT 85.120 66.980 93.160 67.150 ;
        RECT 93.375 65.920 93.545 66.920 ;
        RECT 85.120 65.690 93.160 65.860 ;
        RECT 93.890 65.320 94.060 67.550 ;
        RECT 84.580 65.120 94.060 65.320 ;
        RECT 84.580 62.920 84.750 65.120 ;
        RECT 85.120 64.580 93.160 64.750 ;
        RECT 93.375 63.520 93.545 64.520 ;
        RECT 85.120 63.290 93.160 63.460 ;
        RECT 93.890 62.920 94.060 65.120 ;
        RECT 84.580 62.720 94.060 62.920 ;
        RECT 74.480 62.450 83.810 62.500 ;
        RECT 61.580 57.850 63.480 57.925 ;
        RECT 58.580 57.350 61.180 57.520 ;
        RECT 58.580 48.260 58.750 57.350 ;
        RECT 59.150 48.940 59.320 56.980 ;
        RECT 60.440 48.940 60.610 56.980 ;
        RECT 59.380 48.600 60.380 48.770 ;
        RECT 61.010 48.260 61.180 57.350 ;
        RECT 61.580 48.590 61.750 57.850 ;
        RECT 62.120 57.280 62.580 57.450 ;
        RECT 62.795 49.220 62.965 57.220 ;
        RECT 62.120 48.990 62.580 49.160 ;
        RECT 63.310 48.590 63.480 57.850 ;
        RECT 61.580 48.420 63.480 48.590 ;
        RECT 63.880 57.350 65.730 57.520 ;
        RECT 58.580 48.090 61.180 48.260 ;
        RECT 63.880 48.090 64.050 57.350 ;
        RECT 64.420 56.780 64.880 56.950 ;
        RECT 65.050 48.720 65.220 56.720 ;
        RECT 64.420 48.490 64.880 48.660 ;
        RECT 65.560 48.090 65.730 57.350 ;
        RECT 67.180 55.490 69.280 55.660 ;
        RECT 67.180 50.350 67.350 55.490 ;
        RECT 67.750 51.080 67.920 55.120 ;
        RECT 68.540 51.080 68.710 55.120 ;
        RECT 67.980 50.695 68.480 50.865 ;
        RECT 69.110 50.350 69.280 55.490 ;
        RECT 74.480 53.190 74.650 62.450 ;
        RECT 75.020 61.880 76.060 62.050 ;
        RECT 76.230 53.820 76.400 61.820 ;
        RECT 75.020 53.590 76.060 53.760 ;
        RECT 76.740 53.190 76.950 62.450 ;
        RECT 77.320 61.880 78.360 62.050 ;
        RECT 78.530 53.820 78.700 61.820 ;
        RECT 77.320 53.590 78.360 53.760 ;
        RECT 79.040 53.190 79.250 62.450 ;
        RECT 79.620 61.880 80.660 62.050 ;
        RECT 80.830 53.820 81.000 61.820 ;
        RECT 79.620 53.590 80.660 53.760 ;
        RECT 81.340 53.190 81.550 62.450 ;
        RECT 81.920 61.880 82.960 62.050 ;
        RECT 74.480 53.020 81.550 53.190 ;
        RECT 67.180 50.180 69.280 50.350 ;
        RECT 55.380 47.920 57.810 48.090 ;
        RECT 63.880 47.920 65.730 48.090 ;
        RECT 81.380 48.090 81.550 53.020 ;
        RECT 83.130 48.720 83.300 61.820 ;
        RECT 81.920 48.490 82.960 48.660 ;
        RECT 83.640 48.090 83.810 62.450 ;
        RECT 84.580 60.525 84.750 62.720 ;
        RECT 85.120 62.180 93.160 62.350 ;
        RECT 93.375 61.120 93.545 62.120 ;
        RECT 85.120 60.890 93.160 61.060 ;
        RECT 93.890 60.525 94.060 62.720 ;
        RECT 84.580 60.320 94.060 60.525 ;
        RECT 84.580 58.095 84.750 60.320 ;
        RECT 85.120 59.785 93.160 59.955 ;
        RECT 93.375 58.725 93.545 59.725 ;
        RECT 85.120 58.495 93.160 58.665 ;
        RECT 93.890 58.095 94.060 60.320 ;
        RECT 84.580 57.925 94.060 58.095 ;
        RECT 87.580 57.850 89.480 57.925 ;
        RECT 84.580 57.350 87.180 57.520 ;
        RECT 84.580 48.260 84.750 57.350 ;
        RECT 85.150 48.940 85.320 56.980 ;
        RECT 86.440 48.940 86.610 56.980 ;
        RECT 85.380 48.600 86.380 48.770 ;
        RECT 87.010 48.260 87.180 57.350 ;
        RECT 87.580 48.590 87.750 57.850 ;
        RECT 88.120 57.280 88.580 57.450 ;
        RECT 88.795 49.220 88.965 57.220 ;
        RECT 88.120 48.990 88.580 49.160 ;
        RECT 89.310 48.590 89.480 57.850 ;
        RECT 87.580 48.420 89.480 48.590 ;
        RECT 89.880 57.350 91.730 57.520 ;
        RECT 84.580 48.090 87.180 48.260 ;
        RECT 89.880 48.090 90.050 57.350 ;
        RECT 90.420 56.780 90.880 56.950 ;
        RECT 91.050 48.720 91.220 56.720 ;
        RECT 90.420 48.490 90.880 48.660 ;
        RECT 91.560 48.090 91.730 57.350 ;
        RECT 93.180 55.490 95.280 55.660 ;
        RECT 93.180 50.350 93.350 55.490 ;
        RECT 93.750 51.080 93.920 55.120 ;
        RECT 94.540 51.080 94.710 55.120 ;
        RECT 93.980 50.695 94.480 50.865 ;
        RECT 95.110 50.350 95.280 55.490 ;
        RECT 93.180 50.180 95.280 50.350 ;
        RECT 81.380 47.920 83.810 48.090 ;
        RECT 89.880 47.920 91.730 48.090 ;
        RECT 33.200 46.880 42.800 47.050 ;
        RECT 32.625 46.310 42.300 46.480 ;
        RECT 32.625 44.750 32.870 46.310 ;
        RECT 33.500 45.795 41.500 45.965 ;
        RECT 33.270 45.120 33.440 45.580 ;
        RECT 41.560 45.120 41.730 45.580 ;
        RECT 42.130 44.750 42.300 46.310 ;
        RECT 32.625 44.580 42.300 44.750 ;
        RECT 32.625 41.750 32.795 44.580 ;
        RECT 14.600 41.580 17.200 41.585 ;
        RECT 23.000 41.580 32.795 41.750 ;
        RECT 33.200 44.010 42.630 44.180 ;
        RECT 33.200 41.750 33.370 44.010 ;
        RECT 33.740 43.440 41.780 43.610 ;
        RECT 41.950 42.380 42.120 43.380 ;
        RECT 33.740 42.150 41.780 42.320 ;
        RECT 42.460 41.750 42.630 44.010 ;
        RECT 33.200 41.580 42.630 41.750 ;
        RECT 48.480 42.370 57.910 42.540 ;
        RECT 6.180 40.810 28.220 40.910 ;
        RECT 6.180 40.740 42.800 40.810 ;
        RECT 6.180 31.650 6.350 40.740 ;
        RECT 6.980 40.230 7.980 40.400 ;
        RECT 6.750 32.020 6.920 40.060 ;
        RECT 8.040 32.020 8.210 40.060 ;
        RECT 8.610 31.650 8.780 40.740 ;
        RECT 9.410 40.230 10.410 40.400 ;
        RECT 9.180 32.020 9.350 40.060 ;
        RECT 10.470 32.020 10.640 40.060 ;
        RECT 11.040 31.650 11.210 40.740 ;
        RECT 11.840 40.230 12.840 40.400 ;
        RECT 11.610 32.020 11.780 40.060 ;
        RECT 12.900 32.020 13.070 40.060 ;
        RECT 13.470 31.650 13.640 40.740 ;
        RECT 14.270 40.230 15.270 40.400 ;
        RECT 14.040 32.020 14.210 40.060 ;
        RECT 15.330 32.020 15.500 40.060 ;
        RECT 15.900 31.650 16.070 40.740 ;
        RECT 16.700 40.230 17.700 40.400 ;
        RECT 16.470 32.020 16.640 40.060 ;
        RECT 17.760 32.020 17.930 40.060 ;
        RECT 18.330 31.650 18.500 40.740 ;
        RECT 19.130 40.230 20.130 40.400 ;
        RECT 18.900 32.020 19.070 40.060 ;
        RECT 20.190 32.020 20.360 40.060 ;
        RECT 20.760 31.650 20.930 40.740 ;
        RECT 21.560 40.230 22.560 40.400 ;
        RECT 21.330 32.020 21.500 40.060 ;
        RECT 22.620 32.020 22.790 40.060 ;
        RECT 23.190 31.650 23.360 40.740 ;
        RECT 23.990 40.230 24.990 40.400 ;
        RECT 23.760 32.020 23.930 40.060 ;
        RECT 25.050 32.020 25.220 40.060 ;
        RECT 25.620 31.650 25.790 40.740 ;
        RECT 28.050 40.640 42.800 40.740 ;
        RECT 26.420 40.230 27.420 40.400 ;
        RECT 26.190 32.020 26.360 40.060 ;
        RECT 27.480 32.020 27.650 40.060 ;
        RECT 28.050 38.550 28.270 40.640 ;
        RECT 28.900 40.130 42.000 40.300 ;
        RECT 28.670 38.920 28.840 39.960 ;
        RECT 42.060 38.920 42.230 39.960 ;
        RECT 42.630 38.550 42.800 40.640 ;
        RECT 28.050 38.380 42.800 38.550 ;
        RECT 48.480 40.110 48.650 42.370 ;
        RECT 49.020 41.800 57.060 41.970 ;
        RECT 57.230 40.740 57.400 41.740 ;
        RECT 49.020 40.510 57.060 40.680 ;
        RECT 57.740 40.110 57.910 42.370 ;
        RECT 48.480 39.940 57.910 40.110 ;
        RECT 28.050 38.340 37.700 38.380 ;
        RECT 28.050 36.250 28.270 38.340 ;
        RECT 28.900 37.830 36.900 38.000 ;
        RECT 28.670 36.620 28.840 37.660 ;
        RECT 36.960 36.620 37.130 37.660 ;
        RECT 37.530 36.250 37.700 38.340 ;
        RECT 28.050 36.040 37.700 36.250 ;
        RECT 28.050 33.950 28.270 36.040 ;
        RECT 28.900 35.530 36.900 35.700 ;
        RECT 28.670 34.320 28.840 35.360 ;
        RECT 36.960 34.320 37.130 35.360 ;
        RECT 37.530 33.950 37.700 36.040 ;
        RECT 28.050 33.740 37.700 33.950 ;
        RECT 28.050 31.650 28.270 33.740 ;
        RECT 28.900 33.230 36.900 33.400 ;
        RECT 28.670 32.020 28.840 33.060 ;
        RECT 36.960 32.020 37.130 33.060 ;
        RECT 37.530 31.650 37.700 33.740 ;
        RECT 6.180 31.480 37.700 31.650 ;
        RECT 48.480 37.680 48.650 39.940 ;
        RECT 49.020 39.370 57.060 39.540 ;
        RECT 57.230 38.310 57.400 39.310 ;
        RECT 49.020 38.080 57.060 38.250 ;
        RECT 57.740 37.680 57.910 39.940 ;
        RECT 48.480 37.510 57.910 37.680 ;
        RECT 48.480 35.250 48.650 37.510 ;
        RECT 49.020 36.940 57.060 37.110 ;
        RECT 57.230 35.880 57.400 36.880 ;
        RECT 49.020 35.650 57.060 35.820 ;
        RECT 57.740 35.250 57.910 37.510 ;
        RECT 58.580 42.350 68.060 42.520 ;
        RECT 58.580 40.090 58.750 42.350 ;
        RECT 59.120 41.780 67.160 41.950 ;
        RECT 67.375 40.720 67.545 41.720 ;
        RECT 59.120 40.490 67.160 40.660 ;
        RECT 67.890 40.090 68.060 42.350 ;
        RECT 58.580 39.920 68.060 40.090 ;
        RECT 58.580 37.660 58.750 39.920 ;
        RECT 59.120 39.350 67.160 39.520 ;
        RECT 67.375 38.290 67.545 39.290 ;
        RECT 59.120 38.060 67.160 38.230 ;
        RECT 67.890 37.660 68.060 39.920 ;
        RECT 58.580 37.490 68.060 37.660 ;
        RECT 74.480 42.370 83.910 42.540 ;
        RECT 74.480 40.110 74.650 42.370 ;
        RECT 75.020 41.800 83.060 41.970 ;
        RECT 83.230 40.740 83.400 41.740 ;
        RECT 75.020 40.510 83.060 40.680 ;
        RECT 83.740 40.110 83.910 42.370 ;
        RECT 74.480 39.940 83.910 40.110 ;
        RECT 74.480 37.680 74.650 39.940 ;
        RECT 75.020 39.370 83.060 39.540 ;
        RECT 83.230 38.310 83.400 39.310 ;
        RECT 75.020 38.080 83.060 38.250 ;
        RECT 83.740 37.680 83.910 39.940 ;
        RECT 74.480 37.510 83.910 37.680 ;
        RECT 48.480 35.080 57.910 35.250 ;
        RECT 48.480 32.820 48.650 35.080 ;
        RECT 49.020 34.510 57.060 34.680 ;
        RECT 57.230 33.450 57.400 34.450 ;
        RECT 49.020 33.220 57.060 33.390 ;
        RECT 57.740 32.820 57.910 35.080 ;
        RECT 58.580 36.950 68.010 37.120 ;
        RECT 58.580 34.690 58.750 36.950 ;
        RECT 59.120 36.380 67.160 36.550 ;
        RECT 67.330 35.320 67.500 36.320 ;
        RECT 59.120 35.090 67.160 35.260 ;
        RECT 67.840 34.690 68.010 36.950 ;
        RECT 58.580 34.520 68.010 34.690 ;
        RECT 74.480 35.250 74.650 37.510 ;
        RECT 75.020 36.940 83.060 37.110 ;
        RECT 83.230 35.880 83.400 36.880 ;
        RECT 75.020 35.650 83.060 35.820 ;
        RECT 83.740 35.250 83.910 37.510 ;
        RECT 84.580 42.350 94.060 42.520 ;
        RECT 84.580 40.090 84.750 42.350 ;
        RECT 85.120 41.780 93.160 41.950 ;
        RECT 93.375 40.720 93.545 41.720 ;
        RECT 85.120 40.490 93.160 40.660 ;
        RECT 93.890 40.090 94.060 42.350 ;
        RECT 84.580 39.920 94.060 40.090 ;
        RECT 84.580 37.660 84.750 39.920 ;
        RECT 85.120 39.350 93.160 39.520 ;
        RECT 93.375 38.290 93.545 39.290 ;
        RECT 85.120 38.060 93.160 38.230 ;
        RECT 93.890 37.660 94.060 39.920 ;
        RECT 84.580 37.490 94.060 37.660 ;
        RECT 74.480 35.080 83.910 35.250 ;
        RECT 48.480 32.650 57.910 32.820 ;
        RECT 48.480 30.390 48.650 32.650 ;
        RECT 49.020 32.080 57.060 32.250 ;
        RECT 57.230 31.020 57.400 32.020 ;
        RECT 49.020 30.790 57.060 30.960 ;
        RECT 57.740 30.390 57.910 32.650 ;
        RECT 58.580 33.950 68.060 34.120 ;
        RECT 58.580 31.690 58.750 33.950 ;
        RECT 59.120 33.380 67.160 33.550 ;
        RECT 67.375 32.320 67.545 33.320 ;
        RECT 59.120 32.090 67.160 32.260 ;
        RECT 67.890 31.690 68.060 33.950 ;
        RECT 74.480 32.820 74.650 35.080 ;
        RECT 75.020 34.510 83.060 34.680 ;
        RECT 83.230 33.450 83.400 34.450 ;
        RECT 75.020 33.220 83.060 33.390 ;
        RECT 83.740 32.820 83.910 35.080 ;
        RECT 84.580 36.950 94.010 37.120 ;
        RECT 84.580 34.690 84.750 36.950 ;
        RECT 85.120 36.380 93.160 36.550 ;
        RECT 93.330 35.320 93.500 36.320 ;
        RECT 85.120 35.090 93.160 35.260 ;
        RECT 93.840 34.690 94.010 36.950 ;
        RECT 84.580 34.520 94.010 34.690 ;
        RECT 74.480 32.650 83.910 32.820 ;
        RECT 58.580 31.520 68.065 31.690 ;
        RECT 48.480 30.220 57.910 30.390 ;
        RECT 48.480 27.960 48.650 30.220 ;
        RECT 49.020 29.650 57.060 29.820 ;
        RECT 57.230 28.590 57.400 29.590 ;
        RECT 49.020 28.360 57.060 28.530 ;
        RECT 57.740 27.960 57.910 30.220 ;
        RECT 58.585 29.260 58.755 31.520 ;
        RECT 59.125 30.950 67.165 31.120 ;
        RECT 67.380 29.890 67.550 30.890 ;
        RECT 59.125 29.660 67.165 29.830 ;
        RECT 67.895 29.260 68.065 31.520 ;
        RECT 58.585 29.090 68.065 29.260 ;
        RECT 74.480 30.390 74.650 32.650 ;
        RECT 75.020 32.080 83.060 32.250 ;
        RECT 83.230 31.020 83.400 32.020 ;
        RECT 75.020 30.790 83.060 30.960 ;
        RECT 83.740 30.390 83.910 32.650 ;
        RECT 84.580 33.950 94.060 34.120 ;
        RECT 84.580 31.690 84.750 33.950 ;
        RECT 85.120 33.380 93.160 33.550 ;
        RECT 93.375 32.320 93.545 33.320 ;
        RECT 85.120 32.090 93.160 32.260 ;
        RECT 93.890 31.690 94.060 33.950 ;
        RECT 84.580 31.520 94.065 31.690 ;
        RECT 74.480 30.220 83.910 30.390 ;
        RECT 48.480 27.790 57.910 27.960 ;
        RECT 35.180 26.110 40.660 26.280 ;
        RECT 17.030 25.060 19.630 25.065 ;
        RECT 6.200 24.890 11.230 25.060 ;
        RECT 6.200 15.750 6.370 24.890 ;
        RECT 7.000 24.375 8.000 24.545 ;
        RECT 6.770 16.120 6.940 24.160 ;
        RECT 8.060 16.120 8.230 24.160 ;
        RECT 8.630 15.750 8.800 24.890 ;
        RECT 9.430 24.375 10.430 24.545 ;
        RECT 9.200 16.120 9.370 24.160 ;
        RECT 10.490 16.120 10.660 24.160 ;
        RECT 11.060 15.750 11.230 24.890 ;
        RECT 6.200 15.580 11.230 15.750 ;
        RECT 11.600 24.840 14.200 25.010 ;
        RECT 11.600 15.750 11.770 24.840 ;
        RECT 12.400 24.330 13.400 24.500 ;
        RECT 12.170 16.120 12.340 24.160 ;
        RECT 13.460 16.120 13.630 24.160 ;
        RECT 14.030 15.750 14.200 24.840 ;
        RECT 11.600 15.580 14.200 15.750 ;
        RECT 14.600 24.895 19.630 25.060 ;
        RECT 14.600 24.890 17.200 24.895 ;
        RECT 14.600 15.750 14.770 24.890 ;
        RECT 15.400 24.375 16.400 24.545 ;
        RECT 15.170 16.120 15.340 24.160 ;
        RECT 16.460 16.120 16.630 24.160 ;
        RECT 17.030 15.755 17.200 24.890 ;
        RECT 17.830 24.380 18.830 24.550 ;
        RECT 17.600 16.125 17.770 24.165 ;
        RECT 18.890 16.125 19.060 24.165 ;
        RECT 19.460 15.755 19.630 24.895 ;
        RECT 17.030 15.750 19.630 15.755 ;
        RECT 14.600 15.585 19.630 15.750 ;
        RECT 20.010 24.855 22.610 25.025 ;
        RECT 20.010 15.765 20.180 24.855 ;
        RECT 20.810 24.345 21.810 24.515 ;
        RECT 20.580 16.135 20.750 24.175 ;
        RECT 21.870 16.135 22.040 24.175 ;
        RECT 22.440 15.765 22.610 24.855 ;
        RECT 20.010 15.595 22.610 15.765 ;
        RECT 23.000 24.890 32.795 25.060 ;
        RECT 23.000 15.750 23.170 24.890 ;
        RECT 23.800 24.375 24.800 24.545 ;
        RECT 23.570 16.120 23.740 24.160 ;
        RECT 24.860 16.120 25.030 24.160 ;
        RECT 25.400 15.750 25.600 24.890 ;
        RECT 26.200 24.375 27.200 24.545 ;
        RECT 25.970 16.120 26.140 24.160 ;
        RECT 27.260 16.120 27.430 24.160 ;
        RECT 27.800 15.750 28.000 24.890 ;
        RECT 28.600 24.375 29.600 24.545 ;
        RECT 28.370 16.120 28.540 24.160 ;
        RECT 29.660 16.120 29.830 24.160 ;
        RECT 30.195 15.750 30.400 24.890 ;
        RECT 30.995 24.375 31.995 24.545 ;
        RECT 30.765 16.120 30.935 24.160 ;
        RECT 32.055 16.120 32.225 24.160 ;
        RECT 32.625 20.480 32.795 24.890 ;
        RECT 35.180 24.350 35.350 26.110 ;
        RECT 35.720 25.540 39.760 25.710 ;
        RECT 39.975 24.980 40.145 25.480 ;
        RECT 35.720 24.750 39.760 24.920 ;
        RECT 40.490 24.350 40.660 26.110 ;
        RECT 35.180 24.180 40.660 24.350 ;
        RECT 48.480 25.530 48.650 27.790 ;
        RECT 49.020 27.220 57.060 27.390 ;
        RECT 57.230 26.160 57.400 27.160 ;
        RECT 49.020 25.930 57.060 26.100 ;
        RECT 57.740 25.530 57.910 27.790 ;
        RECT 58.595 28.540 68.025 28.710 ;
        RECT 58.595 26.280 58.765 28.540 ;
        RECT 59.135 27.970 67.175 28.140 ;
        RECT 67.345 26.910 67.515 27.910 ;
        RECT 59.135 26.680 67.175 26.850 ;
        RECT 67.855 26.280 68.025 28.540 ;
        RECT 58.595 26.110 68.025 26.280 ;
        RECT 74.480 27.960 74.650 30.220 ;
        RECT 75.020 29.650 83.060 29.820 ;
        RECT 83.230 28.590 83.400 29.590 ;
        RECT 75.020 28.360 83.060 28.530 ;
        RECT 83.740 27.960 83.910 30.220 ;
        RECT 84.585 29.260 84.755 31.520 ;
        RECT 85.125 30.950 93.165 31.120 ;
        RECT 93.380 29.890 93.550 30.890 ;
        RECT 85.125 29.660 93.165 29.830 ;
        RECT 93.895 29.260 94.065 31.520 ;
        RECT 84.585 29.090 94.065 29.260 ;
        RECT 74.480 27.790 83.910 27.960 ;
        RECT 48.480 25.360 57.910 25.530 ;
        RECT 48.480 23.100 48.650 25.360 ;
        RECT 49.020 24.790 57.060 24.960 ;
        RECT 57.230 23.730 57.400 24.730 ;
        RECT 49.020 23.500 57.060 23.670 ;
        RECT 57.740 23.100 57.910 25.360 ;
        RECT 48.480 22.930 57.910 23.100 ;
        RECT 33.200 22.560 42.800 22.730 ;
        RECT 33.200 21.050 33.370 22.560 ;
        RECT 34.000 22.050 42.000 22.220 ;
        RECT 33.770 21.420 33.940 21.880 ;
        RECT 42.060 21.420 42.230 21.880 ;
        RECT 42.630 21.050 42.800 22.560 ;
        RECT 33.200 20.880 42.800 21.050 ;
        RECT 48.480 20.670 48.650 22.930 ;
        RECT 49.020 22.360 57.060 22.530 ;
        RECT 57.230 21.300 57.400 22.300 ;
        RECT 49.020 21.070 57.060 21.240 ;
        RECT 57.740 20.670 57.910 22.930 ;
        RECT 48.480 20.500 57.910 20.670 ;
        RECT 58.580 25.550 68.060 25.720 ;
        RECT 58.580 23.320 58.750 25.550 ;
        RECT 59.120 24.980 67.160 25.150 ;
        RECT 67.375 23.920 67.545 24.920 ;
        RECT 59.120 23.690 67.160 23.860 ;
        RECT 67.890 23.320 68.060 25.550 ;
        RECT 58.580 23.120 68.060 23.320 ;
        RECT 58.580 20.920 58.750 23.120 ;
        RECT 59.120 22.580 67.160 22.750 ;
        RECT 67.375 21.520 67.545 22.520 ;
        RECT 59.120 21.290 67.160 21.460 ;
        RECT 67.890 20.920 68.060 23.120 ;
        RECT 58.580 20.720 68.060 20.920 ;
        RECT 32.625 20.310 42.300 20.480 ;
        RECT 32.625 18.750 32.870 20.310 ;
        RECT 33.500 19.795 41.500 19.965 ;
        RECT 33.270 19.120 33.440 19.580 ;
        RECT 41.560 19.120 41.730 19.580 ;
        RECT 42.130 18.750 42.300 20.310 ;
        RECT 32.625 18.580 42.300 18.750 ;
        RECT 48.480 20.450 57.810 20.500 ;
        RECT 32.625 15.750 32.795 18.580 ;
        RECT 14.600 15.580 17.200 15.585 ;
        RECT 23.000 15.580 32.795 15.750 ;
        RECT 33.200 18.010 42.630 18.180 ;
        RECT 33.200 15.750 33.370 18.010 ;
        RECT 33.740 17.440 41.780 17.610 ;
        RECT 41.950 16.380 42.120 17.380 ;
        RECT 33.740 16.150 41.780 16.320 ;
        RECT 42.460 15.750 42.630 18.010 ;
        RECT 33.200 15.580 42.630 15.750 ;
        RECT 6.180 14.810 28.220 14.910 ;
        RECT 6.180 14.740 42.800 14.810 ;
        RECT 6.180 5.650 6.350 14.740 ;
        RECT 6.980 14.230 7.980 14.400 ;
        RECT 6.750 6.020 6.920 14.060 ;
        RECT 8.040 6.020 8.210 14.060 ;
        RECT 8.610 5.650 8.780 14.740 ;
        RECT 9.410 14.230 10.410 14.400 ;
        RECT 9.180 6.020 9.350 14.060 ;
        RECT 10.470 6.020 10.640 14.060 ;
        RECT 11.040 5.650 11.210 14.740 ;
        RECT 11.840 14.230 12.840 14.400 ;
        RECT 11.610 6.020 11.780 14.060 ;
        RECT 12.900 6.020 13.070 14.060 ;
        RECT 13.470 5.650 13.640 14.740 ;
        RECT 14.270 14.230 15.270 14.400 ;
        RECT 14.040 6.020 14.210 14.060 ;
        RECT 15.330 6.020 15.500 14.060 ;
        RECT 15.900 5.650 16.070 14.740 ;
        RECT 16.700 14.230 17.700 14.400 ;
        RECT 16.470 6.020 16.640 14.060 ;
        RECT 17.760 6.020 17.930 14.060 ;
        RECT 18.330 5.650 18.500 14.740 ;
        RECT 19.130 14.230 20.130 14.400 ;
        RECT 18.900 6.020 19.070 14.060 ;
        RECT 20.190 6.020 20.360 14.060 ;
        RECT 20.760 5.650 20.930 14.740 ;
        RECT 21.560 14.230 22.560 14.400 ;
        RECT 21.330 6.020 21.500 14.060 ;
        RECT 22.620 6.020 22.790 14.060 ;
        RECT 23.190 5.650 23.360 14.740 ;
        RECT 23.990 14.230 24.990 14.400 ;
        RECT 23.760 6.020 23.930 14.060 ;
        RECT 25.050 6.020 25.220 14.060 ;
        RECT 25.620 5.650 25.790 14.740 ;
        RECT 28.050 14.640 42.800 14.740 ;
        RECT 26.420 14.230 27.420 14.400 ;
        RECT 26.190 6.020 26.360 14.060 ;
        RECT 27.480 6.020 27.650 14.060 ;
        RECT 28.050 12.550 28.270 14.640 ;
        RECT 28.900 14.130 42.000 14.300 ;
        RECT 28.670 12.920 28.840 13.960 ;
        RECT 42.060 12.920 42.230 13.960 ;
        RECT 42.630 12.550 42.800 14.640 ;
        RECT 28.050 12.380 42.800 12.550 ;
        RECT 28.050 12.340 37.700 12.380 ;
        RECT 28.050 10.250 28.270 12.340 ;
        RECT 28.900 11.830 36.900 12.000 ;
        RECT 28.670 10.620 28.840 11.660 ;
        RECT 36.960 10.620 37.130 11.660 ;
        RECT 37.530 10.250 37.700 12.340 ;
        RECT 48.480 11.190 48.650 20.450 ;
        RECT 49.020 19.880 50.060 20.050 ;
        RECT 50.230 11.820 50.400 19.820 ;
        RECT 49.020 11.590 50.060 11.760 ;
        RECT 50.740 11.190 50.950 20.450 ;
        RECT 51.320 19.880 52.360 20.050 ;
        RECT 52.530 11.820 52.700 19.820 ;
        RECT 51.320 11.590 52.360 11.760 ;
        RECT 53.040 11.190 53.250 20.450 ;
        RECT 53.620 19.880 54.660 20.050 ;
        RECT 54.830 11.820 55.000 19.820 ;
        RECT 53.620 11.590 54.660 11.760 ;
        RECT 55.340 11.190 55.550 20.450 ;
        RECT 55.920 19.880 56.960 20.050 ;
        RECT 48.480 11.020 55.550 11.190 ;
        RECT 28.050 10.040 37.700 10.250 ;
        RECT 28.050 7.950 28.270 10.040 ;
        RECT 28.900 9.530 36.900 9.700 ;
        RECT 28.670 8.320 28.840 9.360 ;
        RECT 36.960 8.320 37.130 9.360 ;
        RECT 37.530 7.950 37.700 10.040 ;
        RECT 28.050 7.740 37.700 7.950 ;
        RECT 28.050 5.650 28.270 7.740 ;
        RECT 28.900 7.230 36.900 7.400 ;
        RECT 28.670 6.020 28.840 7.060 ;
        RECT 36.960 6.020 37.130 7.060 ;
        RECT 37.530 5.650 37.700 7.740 ;
        RECT 55.380 6.090 55.550 11.020 ;
        RECT 57.130 6.720 57.300 19.820 ;
        RECT 55.920 6.490 56.960 6.660 ;
        RECT 57.640 6.090 57.810 20.450 ;
        RECT 58.580 18.525 58.750 20.720 ;
        RECT 59.120 20.180 67.160 20.350 ;
        RECT 67.375 19.120 67.545 20.120 ;
        RECT 59.120 18.890 67.160 19.060 ;
        RECT 67.890 18.525 68.060 20.720 ;
        RECT 58.580 18.320 68.060 18.525 ;
        RECT 58.580 16.095 58.750 18.320 ;
        RECT 59.120 17.785 67.160 17.955 ;
        RECT 67.375 16.725 67.545 17.725 ;
        RECT 59.120 16.495 67.160 16.665 ;
        RECT 67.890 16.095 68.060 18.320 ;
        RECT 58.580 15.925 68.060 16.095 ;
        RECT 74.480 25.530 74.650 27.790 ;
        RECT 75.020 27.220 83.060 27.390 ;
        RECT 83.230 26.160 83.400 27.160 ;
        RECT 75.020 25.930 83.060 26.100 ;
        RECT 83.740 25.530 83.910 27.790 ;
        RECT 84.595 28.540 94.025 28.710 ;
        RECT 84.595 26.280 84.765 28.540 ;
        RECT 85.135 27.970 93.175 28.140 ;
        RECT 93.345 26.910 93.515 27.910 ;
        RECT 85.135 26.680 93.175 26.850 ;
        RECT 93.855 26.280 94.025 28.540 ;
        RECT 84.595 26.110 94.025 26.280 ;
        RECT 74.480 25.360 83.910 25.530 ;
        RECT 74.480 23.100 74.650 25.360 ;
        RECT 75.020 24.790 83.060 24.960 ;
        RECT 83.230 23.730 83.400 24.730 ;
        RECT 75.020 23.500 83.060 23.670 ;
        RECT 83.740 23.100 83.910 25.360 ;
        RECT 74.480 22.930 83.910 23.100 ;
        RECT 74.480 20.670 74.650 22.930 ;
        RECT 75.020 22.360 83.060 22.530 ;
        RECT 83.230 21.300 83.400 22.300 ;
        RECT 75.020 21.070 83.060 21.240 ;
        RECT 83.740 20.670 83.910 22.930 ;
        RECT 74.480 20.500 83.910 20.670 ;
        RECT 84.580 25.550 94.060 25.720 ;
        RECT 84.580 23.320 84.750 25.550 ;
        RECT 85.120 24.980 93.160 25.150 ;
        RECT 93.375 23.920 93.545 24.920 ;
        RECT 85.120 23.690 93.160 23.860 ;
        RECT 93.890 23.320 94.060 25.550 ;
        RECT 84.580 23.120 94.060 23.320 ;
        RECT 84.580 20.920 84.750 23.120 ;
        RECT 85.120 22.580 93.160 22.750 ;
        RECT 93.375 21.520 93.545 22.520 ;
        RECT 85.120 21.290 93.160 21.460 ;
        RECT 93.890 20.920 94.060 23.120 ;
        RECT 84.580 20.720 94.060 20.920 ;
        RECT 74.480 20.450 83.810 20.500 ;
        RECT 61.580 15.850 63.480 15.925 ;
        RECT 58.580 15.350 61.180 15.520 ;
        RECT 58.580 6.260 58.750 15.350 ;
        RECT 59.150 6.940 59.320 14.980 ;
        RECT 60.440 6.940 60.610 14.980 ;
        RECT 59.380 6.600 60.380 6.770 ;
        RECT 61.010 6.260 61.180 15.350 ;
        RECT 61.580 6.590 61.750 15.850 ;
        RECT 62.120 15.280 62.580 15.450 ;
        RECT 62.795 7.220 62.965 15.220 ;
        RECT 62.120 6.990 62.580 7.160 ;
        RECT 63.310 6.590 63.480 15.850 ;
        RECT 61.580 6.420 63.480 6.590 ;
        RECT 63.880 15.350 65.730 15.520 ;
        RECT 58.580 6.090 61.180 6.260 ;
        RECT 63.880 6.090 64.050 15.350 ;
        RECT 64.420 14.780 64.880 14.950 ;
        RECT 65.050 6.720 65.220 14.720 ;
        RECT 64.420 6.490 64.880 6.660 ;
        RECT 65.560 6.090 65.730 15.350 ;
        RECT 67.180 13.490 69.280 13.660 ;
        RECT 67.180 8.350 67.350 13.490 ;
        RECT 67.750 9.080 67.920 13.120 ;
        RECT 68.540 9.080 68.710 13.120 ;
        RECT 67.980 8.695 68.480 8.865 ;
        RECT 69.110 8.350 69.280 13.490 ;
        RECT 74.480 11.190 74.650 20.450 ;
        RECT 75.020 19.880 76.060 20.050 ;
        RECT 76.230 11.820 76.400 19.820 ;
        RECT 75.020 11.590 76.060 11.760 ;
        RECT 76.740 11.190 76.950 20.450 ;
        RECT 77.320 19.880 78.360 20.050 ;
        RECT 78.530 11.820 78.700 19.820 ;
        RECT 77.320 11.590 78.360 11.760 ;
        RECT 79.040 11.190 79.250 20.450 ;
        RECT 79.620 19.880 80.660 20.050 ;
        RECT 80.830 11.820 81.000 19.820 ;
        RECT 79.620 11.590 80.660 11.760 ;
        RECT 81.340 11.190 81.550 20.450 ;
        RECT 81.920 19.880 82.960 20.050 ;
        RECT 74.480 11.020 81.550 11.190 ;
        RECT 67.180 8.180 69.280 8.350 ;
        RECT 55.380 5.920 57.810 6.090 ;
        RECT 63.880 5.920 65.730 6.090 ;
        RECT 81.380 6.090 81.550 11.020 ;
        RECT 83.130 6.720 83.300 19.820 ;
        RECT 81.920 6.490 82.960 6.660 ;
        RECT 83.640 6.090 83.810 20.450 ;
        RECT 84.580 18.525 84.750 20.720 ;
        RECT 85.120 20.180 93.160 20.350 ;
        RECT 93.375 19.120 93.545 20.120 ;
        RECT 85.120 18.890 93.160 19.060 ;
        RECT 93.890 18.525 94.060 20.720 ;
        RECT 84.580 18.320 94.060 18.525 ;
        RECT 84.580 16.095 84.750 18.320 ;
        RECT 85.120 17.785 93.160 17.955 ;
        RECT 93.375 16.725 93.545 17.725 ;
        RECT 85.120 16.495 93.160 16.665 ;
        RECT 93.890 16.095 94.060 18.320 ;
        RECT 84.580 15.925 94.060 16.095 ;
        RECT 87.580 15.850 89.480 15.925 ;
        RECT 84.580 15.350 87.180 15.520 ;
        RECT 84.580 6.260 84.750 15.350 ;
        RECT 85.150 6.940 85.320 14.980 ;
        RECT 86.440 6.940 86.610 14.980 ;
        RECT 85.380 6.600 86.380 6.770 ;
        RECT 87.010 6.260 87.180 15.350 ;
        RECT 87.580 6.590 87.750 15.850 ;
        RECT 88.120 15.280 88.580 15.450 ;
        RECT 88.795 7.220 88.965 15.220 ;
        RECT 88.120 6.990 88.580 7.160 ;
        RECT 89.310 6.590 89.480 15.850 ;
        RECT 87.580 6.420 89.480 6.590 ;
        RECT 89.880 15.350 91.730 15.520 ;
        RECT 84.580 6.090 87.180 6.260 ;
        RECT 89.880 6.090 90.050 15.350 ;
        RECT 90.420 14.780 90.880 14.950 ;
        RECT 91.050 6.720 91.220 14.720 ;
        RECT 90.420 6.490 90.880 6.660 ;
        RECT 91.560 6.090 91.730 15.350 ;
        RECT 93.180 13.490 95.280 13.660 ;
        RECT 93.180 8.350 93.350 13.490 ;
        RECT 93.750 9.080 93.920 13.120 ;
        RECT 94.540 9.080 94.710 13.120 ;
        RECT 93.980 8.695 94.480 8.865 ;
        RECT 95.110 8.350 95.280 13.490 ;
        RECT 93.180 8.180 95.280 8.350 ;
        RECT 81.380 5.920 83.810 6.090 ;
        RECT 89.880 5.920 91.730 6.090 ;
        RECT 6.180 5.480 37.700 5.650 ;
      LAYER met1 ;
        RECT 1.000 210.000 99.000 212.000 ;
        RECT 1.000 208.400 3.000 210.000 ;
        RECT 1.000 208.310 36.800 208.400 ;
        RECT 1.000 208.200 39.265 208.310 ;
        RECT 1.000 207.000 3.000 208.200 ;
        RECT 6.220 204.665 6.420 208.200 ;
        RECT 6.720 206.140 6.920 208.200 ;
        RECT 7.220 206.575 7.720 207.300 ;
        RECT 7.220 206.400 7.770 206.575 ;
        RECT 7.230 206.345 7.770 206.400 ;
        RECT 6.720 205.800 6.970 206.140 ;
        RECT 6.170 204.400 6.420 204.665 ;
        RECT 6.170 199.975 6.400 204.400 ;
        RECT 6.740 198.140 6.970 205.800 ;
        RECT 8.030 198.400 8.260 206.140 ;
        RECT 8.620 204.665 8.820 208.200 ;
        RECT 12.120 207.500 12.620 208.000 ;
        RECT 9.720 206.575 10.220 207.300 ;
        RECT 9.660 206.400 10.220 206.575 ;
        RECT 12.120 206.600 12.320 207.500 ;
        RECT 12.120 206.530 12.820 206.600 ;
        RECT 12.120 206.400 13.170 206.530 ;
        RECT 9.660 206.345 10.200 206.400 ;
        RECT 12.120 206.140 12.320 206.400 ;
        RECT 12.630 206.300 13.170 206.400 ;
        RECT 8.600 199.975 8.830 204.665 ;
        RECT 9.170 198.400 9.400 206.140 ;
        RECT 8.030 198.200 9.400 198.400 ;
        RECT 8.030 198.140 8.260 198.200 ;
        RECT 9.170 198.140 9.400 198.200 ;
        RECT 10.460 198.400 10.690 206.140 ;
        RECT 12.120 205.900 12.370 206.140 ;
        RECT 11.570 204.600 11.800 204.630 ;
        RECT 11.570 204.400 11.820 204.600 ;
        RECT 11.570 199.960 11.800 204.400 ;
        RECT 12.140 198.400 12.370 205.900 ;
        RECT 10.460 198.200 12.370 198.400 ;
        RECT 10.460 198.140 10.690 198.200 ;
        RECT 12.140 198.140 12.370 198.200 ;
        RECT 13.430 198.400 13.660 206.140 ;
        RECT 14.520 204.665 14.720 208.200 ;
        RECT 15.120 206.140 15.320 208.200 ;
        RECT 15.620 206.575 16.120 207.300 ;
        RECT 15.620 206.400 16.170 206.575 ;
        RECT 15.630 206.345 16.170 206.400 ;
        RECT 15.120 205.800 15.370 206.140 ;
        RECT 14.520 204.400 14.800 204.665 ;
        RECT 14.570 199.975 14.800 204.400 ;
        RECT 13.430 198.140 13.720 198.400 ;
        RECT 15.140 198.140 15.370 205.800 ;
        RECT 16.430 198.400 16.660 206.140 ;
        RECT 17.020 204.670 17.220 208.200 ;
        RECT 20.820 207.500 21.320 208.000 ;
        RECT 18.020 206.600 18.520 207.300 ;
        RECT 18.020 206.400 20.720 206.600 ;
        RECT 21.020 206.545 21.320 207.500 ;
        RECT 21.020 206.400 21.580 206.545 ;
        RECT 18.060 206.350 18.600 206.400 ;
        RECT 20.520 206.155 20.720 206.400 ;
        RECT 21.040 206.315 21.580 206.400 ;
        RECT 17.000 199.980 17.230 204.670 ;
        RECT 17.570 198.400 17.800 206.145 ;
        RECT 16.430 198.200 17.800 198.400 ;
        RECT 16.430 198.140 16.660 198.200 ;
        RECT 17.570 198.145 17.800 198.200 ;
        RECT 18.860 198.400 19.090 206.145 ;
        RECT 20.520 205.900 20.780 206.155 ;
        RECT 19.980 199.975 20.210 204.645 ;
        RECT 20.550 198.400 20.780 205.900 ;
        RECT 18.860 198.200 20.780 198.400 ;
        RECT 18.860 198.145 19.090 198.200 ;
        RECT 20.550 198.155 20.780 198.200 ;
        RECT 21.840 198.400 22.070 206.155 ;
        RECT 22.920 204.665 23.120 208.200 ;
        RECT 23.520 206.140 23.720 208.200 ;
        RECT 24.020 206.575 24.520 207.300 ;
        RECT 24.020 206.400 24.570 206.575 ;
        RECT 24.030 206.345 24.570 206.400 ;
        RECT 23.520 205.800 23.770 206.140 ;
        RECT 22.920 204.400 23.200 204.665 ;
        RECT 22.970 199.975 23.200 204.400 ;
        RECT 21.840 198.155 22.120 198.400 ;
        RECT 13.520 198.100 13.720 198.140 ;
        RECT 13.520 197.900 14.520 198.100 ;
        RECT 13.620 197.400 14.120 197.700 ;
        RECT 14.320 197.600 14.520 197.900 ;
        RECT 14.320 197.400 16.620 197.600 ;
        RECT 6.620 197.200 14.120 197.400 ;
        RECT 6.620 196.040 6.820 197.200 ;
        RECT 7.220 196.430 7.720 197.000 ;
        RECT 7.210 196.200 7.750 196.430 ;
        RECT 9.120 196.040 9.320 197.200 ;
        RECT 9.620 196.430 10.120 197.000 ;
        RECT 9.620 196.300 10.180 196.430 ;
        RECT 9.640 196.200 10.180 196.300 ;
        RECT 11.520 196.040 11.720 197.200 ;
        RECT 12.020 196.430 12.520 197.000 ;
        RECT 12.020 196.300 12.610 196.430 ;
        RECT 12.070 196.200 12.610 196.300 ;
        RECT 13.920 196.040 14.120 197.200 ;
        RECT 16.420 197.000 16.620 197.400 ;
        RECT 18.520 197.400 19.020 197.700 ;
        RECT 21.920 197.400 22.120 198.155 ;
        RECT 23.540 198.140 23.770 205.800 ;
        RECT 24.830 198.500 25.060 206.140 ;
        RECT 25.320 204.665 25.520 208.200 ;
        RECT 26.420 206.575 26.920 207.300 ;
        RECT 26.420 206.400 26.970 206.575 ;
        RECT 26.430 206.345 26.970 206.400 ;
        RECT 25.320 204.400 25.600 204.665 ;
        RECT 25.370 199.975 25.600 204.400 ;
        RECT 25.940 198.500 26.170 206.140 ;
        RECT 24.830 198.300 26.170 198.500 ;
        RECT 24.830 198.140 25.060 198.300 ;
        RECT 25.940 198.140 26.170 198.300 ;
        RECT 27.230 198.400 27.460 206.140 ;
        RECT 27.720 204.665 27.920 208.200 ;
        RECT 28.320 206.140 28.520 208.200 ;
        RECT 28.820 206.575 29.320 207.300 ;
        RECT 28.820 206.400 29.370 206.575 ;
        RECT 28.830 206.345 29.370 206.400 ;
        RECT 28.320 205.800 28.570 206.140 ;
        RECT 27.720 204.400 28.000 204.665 ;
        RECT 27.770 199.975 28.000 204.400 ;
        RECT 27.230 198.140 27.520 198.400 ;
        RECT 28.340 198.140 28.570 205.800 ;
        RECT 29.630 198.400 29.860 206.140 ;
        RECT 30.120 204.665 30.320 208.200 ;
        RECT 31.920 207.500 32.420 208.000 ;
        RECT 31.220 206.575 31.720 207.300 ;
        RECT 31.220 206.400 31.765 206.575 ;
        RECT 31.225 206.345 31.765 206.400 ;
        RECT 32.120 206.140 32.320 207.500 ;
        RECT 30.120 204.400 30.395 204.665 ;
        RECT 30.165 199.975 30.395 204.400 ;
        RECT 30.735 198.400 30.965 206.140 ;
        RECT 29.630 198.200 30.965 198.400 ;
        RECT 29.630 198.140 29.860 198.200 ;
        RECT 30.735 198.140 30.965 198.200 ;
        RECT 32.025 205.900 32.320 206.140 ;
        RECT 32.025 198.140 32.255 205.900 ;
        RECT 32.620 201.980 32.820 208.200 ;
        RECT 36.575 208.080 39.265 208.200 ;
        RECT 33.400 207.800 33.900 208.000 ;
        RECT 33.400 207.740 36.000 207.800 ;
        RECT 33.400 207.600 39.740 207.740 ;
        RECT 33.400 207.500 33.900 207.600 ;
        RECT 35.740 207.510 39.740 207.600 ;
        RECT 39.945 207.300 40.175 207.460 ;
        RECT 40.900 207.300 41.600 207.800 ;
        RECT 33.420 206.800 33.920 207.300 ;
        RECT 39.945 207.100 41.600 207.300 ;
        RECT 41.900 207.100 42.600 207.800 ;
        RECT 39.945 207.000 40.175 207.100 ;
        RECT 33.170 203.700 33.400 204.245 ;
        RECT 33.120 203.365 33.400 203.700 ;
        RECT 33.720 203.860 33.920 206.800 ;
        RECT 35.740 206.800 39.740 206.950 ;
        RECT 35.740 206.720 44.100 206.800 ;
        RECT 39.400 206.600 44.100 206.720 ;
        RECT 38.020 204.500 38.520 205.000 ;
        RECT 38.020 204.250 38.220 204.500 ;
        RECT 35.980 204.020 40.020 204.250 ;
        RECT 33.720 203.600 33.970 203.860 ;
        RECT 42.030 203.700 42.260 203.860 ;
        RECT 33.740 203.440 33.970 203.600 ;
        RECT 42.020 203.440 42.260 203.700 ;
        RECT 33.120 202.900 33.320 203.365 ;
        RECT 42.020 202.900 42.220 203.440 ;
        RECT 33.120 202.700 43.720 202.900 ;
        RECT 39.220 201.995 43.320 202.000 ;
        RECT 32.620 201.500 32.900 201.980 ;
        RECT 35.480 201.800 43.320 201.995 ;
        RECT 35.480 201.765 39.520 201.800 ;
        RECT 33.240 201.500 33.470 201.560 ;
        RECT 32.620 201.300 33.470 201.500 ;
        RECT 41.530 201.400 41.760 201.560 ;
        RECT 32.670 201.080 32.900 201.300 ;
        RECT 33.240 201.140 33.470 201.300 ;
        RECT 41.520 201.200 42.920 201.400 ;
        RECT 41.530 201.140 41.760 201.200 ;
        RECT 42.720 200.000 42.920 201.200 ;
        RECT 42.420 199.700 42.920 200.000 ;
        RECT 41.420 199.640 42.920 199.700 ;
        RECT 33.760 199.500 42.920 199.640 ;
        RECT 33.760 199.410 41.760 199.500 ;
        RECT 33.170 198.800 33.400 199.280 ;
        RECT 41.920 199.100 42.150 199.150 ;
        RECT 43.120 199.100 43.320 201.800 ;
        RECT 41.920 198.900 43.320 199.100 ;
        RECT 33.170 198.480 33.420 198.800 ;
        RECT 41.920 198.610 42.150 198.900 ;
        RECT 42.420 198.600 42.920 198.900 ;
        RECT 27.320 197.400 27.520 198.140 ;
        RECT 33.220 197.800 33.420 198.480 ;
        RECT 33.760 198.120 41.760 198.350 ;
        RECT 33.820 197.800 34.020 198.120 ;
        RECT 43.520 197.800 43.720 202.700 ;
        RECT 33.220 197.600 43.720 197.800 ;
        RECT 18.520 197.200 26.320 197.400 ;
        RECT 27.320 197.200 42.220 197.400 ;
        RECT 14.520 196.430 15.020 197.000 ;
        RECT 16.420 196.800 17.420 197.000 ;
        RECT 14.500 196.200 15.040 196.430 ;
        RECT 16.420 196.040 16.620 196.800 ;
        RECT 16.920 196.430 17.420 196.800 ;
        RECT 16.920 196.300 17.470 196.430 ;
        RECT 16.930 196.200 17.470 196.300 ;
        RECT 18.820 196.040 19.020 197.200 ;
        RECT 19.420 196.430 19.920 197.000 ;
        RECT 19.360 196.300 19.920 196.430 ;
        RECT 19.360 196.200 19.900 196.300 ;
        RECT 21.220 196.040 21.420 197.200 ;
        RECT 21.820 196.430 22.320 197.000 ;
        RECT 21.790 196.200 22.330 196.430 ;
        RECT 23.720 196.040 23.920 197.200 ;
        RECT 24.220 196.430 24.720 197.000 ;
        RECT 24.220 196.200 24.760 196.430 ;
        RECT 26.120 196.040 26.320 197.200 ;
        RECT 26.620 196.430 27.120 197.000 ;
        RECT 26.620 196.300 27.190 196.430 ;
        RECT 26.650 196.200 27.190 196.300 ;
        RECT 32.155 196.300 38.745 196.330 ;
        RECT 42.020 196.300 42.220 197.200 ;
        RECT 32.155 196.100 42.220 196.300 ;
        RECT 6.620 195.800 6.950 196.040 ;
        RECT 6.720 188.040 6.950 195.800 ;
        RECT 8.010 188.300 8.240 196.040 ;
        RECT 9.120 195.800 9.380 196.040 ;
        RECT 8.010 188.040 8.320 188.300 ;
        RECT 9.150 188.040 9.380 195.800 ;
        RECT 10.440 188.300 10.670 196.040 ;
        RECT 11.520 195.800 11.810 196.040 ;
        RECT 10.440 188.040 10.720 188.300 ;
        RECT 11.580 188.040 11.810 195.800 ;
        RECT 12.870 188.300 13.100 196.040 ;
        RECT 13.920 195.800 14.240 196.040 ;
        RECT 12.870 188.040 13.120 188.300 ;
        RECT 14.010 188.040 14.240 195.800 ;
        RECT 15.300 188.300 15.530 196.040 ;
        RECT 16.420 195.800 16.670 196.040 ;
        RECT 15.300 188.040 15.620 188.300 ;
        RECT 16.440 188.040 16.670 195.800 ;
        RECT 17.730 188.300 17.960 196.040 ;
        RECT 18.820 195.800 19.100 196.040 ;
        RECT 17.730 188.040 18.020 188.300 ;
        RECT 18.870 188.040 19.100 195.800 ;
        RECT 20.160 188.300 20.390 196.040 ;
        RECT 21.220 195.800 21.530 196.040 ;
        RECT 20.160 188.040 20.420 188.300 ;
        RECT 21.300 188.040 21.530 195.800 ;
        RECT 22.590 188.040 22.820 196.040 ;
        RECT 23.720 195.800 23.960 196.040 ;
        RECT 23.730 188.040 23.960 195.800 ;
        RECT 25.020 188.300 25.250 196.040 ;
        RECT 26.120 195.800 26.390 196.040 ;
        RECT 25.020 188.040 25.320 188.300 ;
        RECT 26.160 188.040 26.390 195.800 ;
        RECT 27.450 188.300 27.680 196.040 ;
        RECT 42.020 195.940 42.220 196.100 ;
        RECT 28.640 195.200 28.870 195.940 ;
        RECT 42.020 195.600 42.260 195.940 ;
        RECT 28.620 194.940 28.870 195.200 ;
        RECT 42.030 195.200 42.260 195.600 ;
        RECT 42.520 195.200 43.020 195.500 ;
        RECT 42.030 195.000 43.020 195.200 ;
        RECT 42.030 194.940 42.260 195.000 ;
        RECT 28.620 193.640 28.820 194.940 ;
        RECT 31.800 194.350 39.100 194.580 ;
        RECT 30.880 194.000 34.920 194.030 ;
        RECT 38.120 194.000 38.620 194.200 ;
        RECT 30.880 193.800 38.620 194.000 ;
        RECT 38.120 193.700 38.620 193.800 ;
        RECT 38.820 193.800 39.020 194.350 ;
        RECT 43.220 193.800 43.420 197.600 ;
        RECT 28.620 193.300 28.870 193.640 ;
        RECT 28.640 192.640 28.870 193.300 ;
        RECT 36.930 193.000 37.160 193.640 ;
        RECT 38.820 193.600 43.420 193.800 ;
        RECT 37.420 193.000 37.920 193.200 ;
        RECT 36.930 192.700 37.920 193.000 ;
        RECT 36.930 192.640 37.160 192.700 ;
        RECT 38.820 192.500 39.020 193.600 ;
        RECT 37.420 192.300 39.020 192.500 ;
        RECT 35.020 192.280 37.620 192.300 ;
        RECT 30.525 192.200 37.620 192.280 ;
        RECT 28.020 192.100 37.620 192.200 ;
        RECT 28.020 192.050 35.275 192.100 ;
        RECT 28.020 192.000 30.820 192.050 ;
        RECT 28.020 189.900 28.220 192.000 ;
        RECT 30.880 191.700 34.920 191.730 ;
        RECT 38.120 191.700 38.620 192.000 ;
        RECT 30.880 191.500 38.620 191.700 ;
        RECT 28.640 190.700 28.870 191.340 ;
        RECT 28.620 190.340 28.870 190.700 ;
        RECT 36.930 190.700 37.160 191.340 ;
        RECT 37.420 190.700 37.920 190.900 ;
        RECT 36.930 190.400 37.920 190.700 ;
        RECT 36.930 190.340 37.160 190.400 ;
        RECT 28.620 189.900 28.820 190.340 ;
        RECT 30.525 189.900 35.275 189.980 ;
        RECT 28.020 189.750 35.275 189.900 ;
        RECT 28.020 189.700 30.820 189.750 ;
        RECT 27.450 188.040 27.720 188.300 ;
        RECT 6.220 187.600 6.720 187.900 ;
        RECT 7.080 187.600 7.880 187.680 ;
        RECT 6.220 187.450 7.880 187.600 ;
        RECT 6.220 187.400 7.220 187.450 ;
        RECT 8.120 187.200 8.320 188.040 ;
        RECT 8.720 187.600 9.220 187.900 ;
        RECT 9.510 187.600 10.310 187.680 ;
        RECT 8.720 187.450 10.310 187.600 ;
        RECT 8.720 187.400 9.720 187.450 ;
        RECT 10.520 187.200 10.720 188.040 ;
        RECT 11.120 187.600 11.620 187.900 ;
        RECT 11.940 187.600 12.740 187.680 ;
        RECT 11.120 187.450 12.740 187.600 ;
        RECT 11.120 187.400 12.120 187.450 ;
        RECT 12.920 187.200 13.120 188.040 ;
        RECT 13.520 187.600 14.020 187.900 ;
        RECT 14.370 187.600 15.170 187.680 ;
        RECT 13.520 187.450 15.170 187.600 ;
        RECT 13.520 187.400 14.620 187.450 ;
        RECT 15.420 187.200 15.620 188.040 ;
        RECT 15.920 187.600 16.420 187.900 ;
        RECT 16.800 187.600 17.600 187.680 ;
        RECT 17.820 187.600 18.020 188.040 ;
        RECT 15.920 187.400 18.020 187.600 ;
        RECT 18.420 187.600 18.920 187.900 ;
        RECT 19.230 187.600 20.030 187.680 ;
        RECT 18.420 187.450 20.030 187.600 ;
        RECT 18.420 187.400 19.420 187.450 ;
        RECT 20.220 187.200 20.420 188.040 ;
        RECT 20.820 187.600 21.320 187.900 ;
        RECT 21.660 187.600 22.460 187.680 ;
        RECT 20.820 187.450 22.460 187.600 ;
        RECT 20.820 187.400 21.820 187.450 ;
        RECT 22.620 187.200 22.820 188.040 ;
        RECT 23.320 187.600 23.820 187.900 ;
        RECT 24.090 187.600 24.890 187.680 ;
        RECT 23.320 187.450 24.890 187.600 ;
        RECT 23.320 187.400 24.320 187.450 ;
        RECT 25.120 187.200 25.320 188.040 ;
        RECT 25.720 187.600 26.220 187.900 ;
        RECT 26.520 187.600 27.320 187.680 ;
        RECT 25.720 187.450 27.320 187.600 ;
        RECT 25.720 187.400 26.820 187.450 ;
        RECT 27.520 187.200 27.720 188.040 ;
        RECT 28.020 187.900 28.220 189.700 ;
        RECT 30.880 189.400 34.920 189.430 ;
        RECT 38.120 189.400 38.620 189.700 ;
        RECT 30.880 189.200 38.620 189.400 ;
        RECT 28.640 188.400 28.870 189.040 ;
        RECT 28.620 188.040 28.870 188.400 ;
        RECT 36.930 188.300 37.160 189.040 ;
        RECT 37.420 188.300 37.920 188.500 ;
        RECT 36.930 188.040 37.920 188.300 ;
        RECT 28.620 187.900 28.820 188.040 ;
        RECT 28.020 187.600 28.820 187.900 ;
        RECT 37.020 188.000 37.920 188.040 ;
        RECT 30.525 187.600 35.275 187.680 ;
        RECT 28.020 187.450 35.275 187.600 ;
        RECT 28.020 187.400 30.820 187.450 ;
        RECT 37.020 187.200 37.220 188.000 ;
        RECT 8.120 187.000 37.220 187.200 ;
        RECT 2.300 182.310 36.900 182.400 ;
        RECT 2.300 182.200 39.265 182.310 ;
        RECT 2.300 181.700 3.000 182.200 ;
        RECT 6.220 178.665 6.420 182.200 ;
        RECT 6.720 180.140 6.920 182.200 ;
        RECT 7.220 180.575 7.720 181.300 ;
        RECT 7.220 180.400 7.770 180.575 ;
        RECT 7.230 180.345 7.770 180.400 ;
        RECT 6.720 179.800 6.970 180.140 ;
        RECT 6.170 178.400 6.420 178.665 ;
        RECT 6.170 173.975 6.400 178.400 ;
        RECT 6.740 172.140 6.970 179.800 ;
        RECT 8.030 172.400 8.260 180.140 ;
        RECT 8.620 178.665 8.820 182.200 ;
        RECT 12.120 181.500 12.620 182.000 ;
        RECT 9.720 180.575 10.220 181.300 ;
        RECT 9.660 180.400 10.220 180.575 ;
        RECT 12.120 180.600 12.320 181.500 ;
        RECT 12.120 180.530 12.820 180.600 ;
        RECT 12.120 180.400 13.170 180.530 ;
        RECT 9.660 180.345 10.200 180.400 ;
        RECT 12.120 180.140 12.320 180.400 ;
        RECT 12.630 180.300 13.170 180.400 ;
        RECT 8.600 173.975 8.830 178.665 ;
        RECT 9.170 172.400 9.400 180.140 ;
        RECT 8.030 172.200 9.400 172.400 ;
        RECT 8.030 172.140 8.260 172.200 ;
        RECT 9.170 172.140 9.400 172.200 ;
        RECT 10.460 172.400 10.690 180.140 ;
        RECT 12.120 179.900 12.370 180.140 ;
        RECT 11.570 178.600 11.800 178.630 ;
        RECT 11.570 178.400 11.820 178.600 ;
        RECT 11.570 173.960 11.800 178.400 ;
        RECT 12.140 172.400 12.370 179.900 ;
        RECT 10.460 172.200 12.370 172.400 ;
        RECT 10.460 172.140 10.690 172.200 ;
        RECT 12.140 172.140 12.370 172.200 ;
        RECT 13.430 172.400 13.660 180.140 ;
        RECT 14.520 178.665 14.720 182.200 ;
        RECT 15.120 180.140 15.320 182.200 ;
        RECT 15.620 180.575 16.120 181.300 ;
        RECT 15.620 180.400 16.170 180.575 ;
        RECT 15.630 180.345 16.170 180.400 ;
        RECT 15.120 179.800 15.370 180.140 ;
        RECT 14.520 178.400 14.800 178.665 ;
        RECT 14.570 173.975 14.800 178.400 ;
        RECT 13.430 172.140 13.720 172.400 ;
        RECT 15.140 172.140 15.370 179.800 ;
        RECT 16.430 172.400 16.660 180.140 ;
        RECT 17.020 178.670 17.220 182.200 ;
        RECT 20.820 181.500 21.320 182.000 ;
        RECT 18.020 180.600 18.520 181.300 ;
        RECT 18.020 180.400 20.720 180.600 ;
        RECT 21.020 180.545 21.320 181.500 ;
        RECT 21.020 180.400 21.580 180.545 ;
        RECT 18.060 180.350 18.600 180.400 ;
        RECT 20.520 180.155 20.720 180.400 ;
        RECT 21.040 180.315 21.580 180.400 ;
        RECT 17.000 173.980 17.230 178.670 ;
        RECT 17.570 172.400 17.800 180.145 ;
        RECT 16.430 172.200 17.800 172.400 ;
        RECT 16.430 172.140 16.660 172.200 ;
        RECT 17.570 172.145 17.800 172.200 ;
        RECT 18.860 172.400 19.090 180.145 ;
        RECT 20.520 179.900 20.780 180.155 ;
        RECT 19.980 173.975 20.210 178.645 ;
        RECT 20.550 172.400 20.780 179.900 ;
        RECT 18.860 172.200 20.780 172.400 ;
        RECT 18.860 172.145 19.090 172.200 ;
        RECT 20.550 172.155 20.780 172.200 ;
        RECT 21.840 172.400 22.070 180.155 ;
        RECT 22.920 178.665 23.120 182.200 ;
        RECT 23.520 180.140 23.720 182.200 ;
        RECT 24.020 180.575 24.520 181.300 ;
        RECT 24.020 180.400 24.570 180.575 ;
        RECT 24.030 180.345 24.570 180.400 ;
        RECT 23.520 179.800 23.770 180.140 ;
        RECT 22.920 178.400 23.200 178.665 ;
        RECT 22.970 173.975 23.200 178.400 ;
        RECT 21.840 172.155 22.120 172.400 ;
        RECT 13.520 172.100 13.720 172.140 ;
        RECT 13.520 171.900 14.520 172.100 ;
        RECT 13.620 171.400 14.120 171.700 ;
        RECT 14.320 171.600 14.520 171.900 ;
        RECT 14.320 171.400 16.620 171.600 ;
        RECT 6.620 171.200 14.120 171.400 ;
        RECT 6.620 170.040 6.820 171.200 ;
        RECT 7.220 170.430 7.720 171.000 ;
        RECT 7.210 170.200 7.750 170.430 ;
        RECT 9.120 170.040 9.320 171.200 ;
        RECT 9.620 170.430 10.120 171.000 ;
        RECT 9.620 170.300 10.180 170.430 ;
        RECT 9.640 170.200 10.180 170.300 ;
        RECT 11.520 170.040 11.720 171.200 ;
        RECT 12.020 170.430 12.520 171.000 ;
        RECT 12.020 170.300 12.610 170.430 ;
        RECT 12.070 170.200 12.610 170.300 ;
        RECT 13.920 170.040 14.120 171.200 ;
        RECT 16.420 171.000 16.620 171.400 ;
        RECT 18.520 171.400 19.020 171.700 ;
        RECT 21.920 171.400 22.120 172.155 ;
        RECT 23.540 172.140 23.770 179.800 ;
        RECT 24.830 172.500 25.060 180.140 ;
        RECT 25.320 178.665 25.520 182.200 ;
        RECT 26.420 180.575 26.920 181.300 ;
        RECT 26.420 180.400 26.970 180.575 ;
        RECT 26.430 180.345 26.970 180.400 ;
        RECT 25.320 178.400 25.600 178.665 ;
        RECT 25.370 173.975 25.600 178.400 ;
        RECT 25.940 172.500 26.170 180.140 ;
        RECT 24.830 172.300 26.170 172.500 ;
        RECT 24.830 172.140 25.060 172.300 ;
        RECT 25.940 172.140 26.170 172.300 ;
        RECT 27.230 172.400 27.460 180.140 ;
        RECT 27.720 178.665 27.920 182.200 ;
        RECT 28.320 180.140 28.520 182.200 ;
        RECT 28.820 180.575 29.320 181.300 ;
        RECT 28.820 180.400 29.370 180.575 ;
        RECT 28.830 180.345 29.370 180.400 ;
        RECT 28.320 179.800 28.570 180.140 ;
        RECT 27.720 178.400 28.000 178.665 ;
        RECT 27.770 173.975 28.000 178.400 ;
        RECT 27.230 172.140 27.520 172.400 ;
        RECT 28.340 172.140 28.570 179.800 ;
        RECT 29.630 172.400 29.860 180.140 ;
        RECT 30.120 178.665 30.320 182.200 ;
        RECT 31.920 181.500 32.420 182.000 ;
        RECT 31.220 180.575 31.720 181.300 ;
        RECT 31.220 180.400 31.765 180.575 ;
        RECT 31.225 180.345 31.765 180.400 ;
        RECT 32.120 180.140 32.320 181.500 ;
        RECT 30.120 178.400 30.395 178.665 ;
        RECT 30.165 173.975 30.395 178.400 ;
        RECT 30.735 172.400 30.965 180.140 ;
        RECT 29.630 172.200 30.965 172.400 ;
        RECT 29.630 172.140 29.860 172.200 ;
        RECT 30.735 172.140 30.965 172.200 ;
        RECT 32.025 179.900 32.320 180.140 ;
        RECT 32.025 172.140 32.255 179.900 ;
        RECT 32.620 175.980 32.820 182.200 ;
        RECT 36.575 182.080 39.265 182.200 ;
        RECT 33.400 181.800 33.900 182.000 ;
        RECT 33.400 181.740 36.000 181.800 ;
        RECT 33.400 181.600 39.740 181.740 ;
        RECT 33.400 181.500 33.900 181.600 ;
        RECT 35.740 181.510 39.740 181.600 ;
        RECT 39.945 181.300 40.175 181.460 ;
        RECT 40.900 181.300 41.600 181.800 ;
        RECT 33.420 180.800 33.920 181.300 ;
        RECT 39.945 181.100 41.600 181.300 ;
        RECT 41.900 181.100 42.600 181.800 ;
        RECT 39.945 181.000 40.175 181.100 ;
        RECT 33.170 177.700 33.400 178.245 ;
        RECT 33.120 177.365 33.400 177.700 ;
        RECT 33.720 177.860 33.920 180.800 ;
        RECT 35.740 180.800 39.740 180.950 ;
        RECT 43.900 180.800 44.100 206.600 ;
        RECT 35.740 180.720 44.100 180.800 ;
        RECT 39.400 180.600 44.100 180.720 ;
        RECT 38.020 178.500 38.520 179.000 ;
        RECT 38.020 178.250 38.220 178.500 ;
        RECT 35.980 178.020 40.020 178.250 ;
        RECT 33.720 177.600 33.970 177.860 ;
        RECT 42.030 177.700 42.260 177.860 ;
        RECT 33.740 177.440 33.970 177.600 ;
        RECT 42.020 177.440 42.260 177.700 ;
        RECT 33.120 176.900 33.320 177.365 ;
        RECT 42.020 176.900 42.220 177.440 ;
        RECT 33.120 176.700 43.720 176.900 ;
        RECT 39.220 175.995 43.320 176.000 ;
        RECT 32.620 175.500 32.900 175.980 ;
        RECT 35.480 175.800 43.320 175.995 ;
        RECT 35.480 175.765 39.520 175.800 ;
        RECT 33.240 175.500 33.470 175.560 ;
        RECT 32.620 175.300 33.470 175.500 ;
        RECT 41.530 175.400 41.760 175.560 ;
        RECT 32.670 175.080 32.900 175.300 ;
        RECT 33.240 175.140 33.470 175.300 ;
        RECT 41.520 175.200 42.920 175.400 ;
        RECT 41.530 175.140 41.760 175.200 ;
        RECT 42.720 174.000 42.920 175.200 ;
        RECT 42.420 173.700 42.920 174.000 ;
        RECT 41.420 173.640 42.920 173.700 ;
        RECT 33.760 173.500 42.920 173.640 ;
        RECT 33.760 173.410 41.760 173.500 ;
        RECT 33.170 172.800 33.400 173.280 ;
        RECT 41.920 173.100 42.150 173.150 ;
        RECT 43.120 173.100 43.320 175.800 ;
        RECT 41.920 172.900 43.320 173.100 ;
        RECT 33.170 172.480 33.420 172.800 ;
        RECT 41.920 172.610 42.150 172.900 ;
        RECT 42.420 172.600 42.920 172.900 ;
        RECT 27.320 171.400 27.520 172.140 ;
        RECT 33.220 171.800 33.420 172.480 ;
        RECT 33.760 172.120 41.760 172.350 ;
        RECT 33.820 171.800 34.020 172.120 ;
        RECT 43.520 171.800 43.720 176.700 ;
        RECT 33.220 171.600 43.720 171.800 ;
        RECT 18.520 171.200 26.320 171.400 ;
        RECT 27.320 171.200 42.220 171.400 ;
        RECT 14.520 170.430 15.020 171.000 ;
        RECT 16.420 170.800 17.420 171.000 ;
        RECT 14.500 170.200 15.040 170.430 ;
        RECT 16.420 170.040 16.620 170.800 ;
        RECT 16.920 170.430 17.420 170.800 ;
        RECT 16.920 170.300 17.470 170.430 ;
        RECT 16.930 170.200 17.470 170.300 ;
        RECT 18.820 170.040 19.020 171.200 ;
        RECT 19.420 170.430 19.920 171.000 ;
        RECT 19.360 170.300 19.920 170.430 ;
        RECT 19.360 170.200 19.900 170.300 ;
        RECT 21.220 170.040 21.420 171.200 ;
        RECT 21.820 170.430 22.320 171.000 ;
        RECT 21.790 170.200 22.330 170.430 ;
        RECT 23.720 170.040 23.920 171.200 ;
        RECT 24.220 170.430 24.720 171.000 ;
        RECT 24.220 170.200 24.760 170.430 ;
        RECT 26.120 170.040 26.320 171.200 ;
        RECT 26.620 170.430 27.120 171.000 ;
        RECT 26.620 170.300 27.190 170.430 ;
        RECT 26.650 170.200 27.190 170.300 ;
        RECT 32.155 170.300 38.745 170.330 ;
        RECT 42.020 170.300 42.220 171.200 ;
        RECT 32.155 170.100 42.220 170.300 ;
        RECT 6.620 169.800 6.950 170.040 ;
        RECT 6.720 162.040 6.950 169.800 ;
        RECT 8.010 162.300 8.240 170.040 ;
        RECT 9.120 169.800 9.380 170.040 ;
        RECT 8.010 162.040 8.320 162.300 ;
        RECT 9.150 162.040 9.380 169.800 ;
        RECT 10.440 162.300 10.670 170.040 ;
        RECT 11.520 169.800 11.810 170.040 ;
        RECT 10.440 162.040 10.720 162.300 ;
        RECT 11.580 162.040 11.810 169.800 ;
        RECT 12.870 162.300 13.100 170.040 ;
        RECT 13.920 169.800 14.240 170.040 ;
        RECT 12.870 162.040 13.120 162.300 ;
        RECT 14.010 162.040 14.240 169.800 ;
        RECT 15.300 162.300 15.530 170.040 ;
        RECT 16.420 169.800 16.670 170.040 ;
        RECT 15.300 162.040 15.620 162.300 ;
        RECT 16.440 162.040 16.670 169.800 ;
        RECT 17.730 162.300 17.960 170.040 ;
        RECT 18.820 169.800 19.100 170.040 ;
        RECT 17.730 162.040 18.020 162.300 ;
        RECT 18.870 162.040 19.100 169.800 ;
        RECT 20.160 162.300 20.390 170.040 ;
        RECT 21.220 169.800 21.530 170.040 ;
        RECT 20.160 162.040 20.420 162.300 ;
        RECT 21.300 162.040 21.530 169.800 ;
        RECT 22.590 162.040 22.820 170.040 ;
        RECT 23.720 169.800 23.960 170.040 ;
        RECT 23.730 162.040 23.960 169.800 ;
        RECT 25.020 162.300 25.250 170.040 ;
        RECT 26.120 169.800 26.390 170.040 ;
        RECT 25.020 162.040 25.320 162.300 ;
        RECT 26.160 162.040 26.390 169.800 ;
        RECT 27.450 162.300 27.680 170.040 ;
        RECT 42.020 169.940 42.220 170.100 ;
        RECT 28.640 169.200 28.870 169.940 ;
        RECT 42.020 169.600 42.260 169.940 ;
        RECT 28.620 168.940 28.870 169.200 ;
        RECT 42.030 169.200 42.260 169.600 ;
        RECT 42.520 169.200 43.020 169.500 ;
        RECT 42.030 169.000 43.020 169.200 ;
        RECT 42.030 168.940 42.260 169.000 ;
        RECT 28.620 167.640 28.820 168.940 ;
        RECT 31.800 168.350 39.100 168.580 ;
        RECT 30.880 168.000 34.920 168.030 ;
        RECT 38.120 168.000 38.620 168.200 ;
        RECT 30.880 167.800 38.620 168.000 ;
        RECT 38.120 167.700 38.620 167.800 ;
        RECT 38.820 167.800 39.020 168.350 ;
        RECT 43.220 167.800 43.420 171.600 ;
        RECT 28.620 167.300 28.870 167.640 ;
        RECT 28.640 166.640 28.870 167.300 ;
        RECT 36.930 167.000 37.160 167.640 ;
        RECT 38.820 167.600 43.420 167.800 ;
        RECT 37.420 167.000 37.920 167.200 ;
        RECT 36.930 166.700 37.920 167.000 ;
        RECT 36.930 166.640 37.160 166.700 ;
        RECT 38.820 166.500 39.020 167.600 ;
        RECT 37.420 166.300 39.020 166.500 ;
        RECT 35.020 166.280 37.620 166.300 ;
        RECT 30.525 166.200 37.620 166.280 ;
        RECT 28.020 166.100 37.620 166.200 ;
        RECT 28.020 166.050 35.275 166.100 ;
        RECT 28.020 166.000 30.820 166.050 ;
        RECT 28.020 163.900 28.220 166.000 ;
        RECT 30.880 165.700 34.920 165.730 ;
        RECT 38.120 165.700 38.620 166.000 ;
        RECT 30.880 165.500 38.620 165.700 ;
        RECT 28.640 164.700 28.870 165.340 ;
        RECT 28.620 164.340 28.870 164.700 ;
        RECT 36.930 164.700 37.160 165.340 ;
        RECT 37.420 164.700 37.920 164.900 ;
        RECT 36.930 164.400 37.920 164.700 ;
        RECT 36.930 164.340 37.160 164.400 ;
        RECT 28.620 163.900 28.820 164.340 ;
        RECT 30.525 163.900 35.275 163.980 ;
        RECT 28.020 163.750 35.275 163.900 ;
        RECT 28.020 163.700 30.820 163.750 ;
        RECT 27.450 162.040 27.720 162.300 ;
        RECT 6.220 161.600 6.720 161.900 ;
        RECT 7.080 161.600 7.880 161.680 ;
        RECT 6.220 161.450 7.880 161.600 ;
        RECT 6.220 161.400 7.220 161.450 ;
        RECT 8.120 161.200 8.320 162.040 ;
        RECT 8.720 161.600 9.220 161.900 ;
        RECT 9.510 161.600 10.310 161.680 ;
        RECT 8.720 161.450 10.310 161.600 ;
        RECT 8.720 161.400 9.720 161.450 ;
        RECT 10.520 161.200 10.720 162.040 ;
        RECT 11.120 161.600 11.620 161.900 ;
        RECT 11.940 161.600 12.740 161.680 ;
        RECT 11.120 161.450 12.740 161.600 ;
        RECT 11.120 161.400 12.120 161.450 ;
        RECT 12.920 161.200 13.120 162.040 ;
        RECT 13.520 161.600 14.020 161.900 ;
        RECT 14.370 161.600 15.170 161.680 ;
        RECT 13.520 161.450 15.170 161.600 ;
        RECT 13.520 161.400 14.620 161.450 ;
        RECT 15.420 161.200 15.620 162.040 ;
        RECT 15.920 161.600 16.420 161.900 ;
        RECT 16.800 161.600 17.600 161.680 ;
        RECT 17.820 161.600 18.020 162.040 ;
        RECT 15.920 161.400 18.020 161.600 ;
        RECT 18.420 161.600 18.920 161.900 ;
        RECT 19.230 161.600 20.030 161.680 ;
        RECT 18.420 161.450 20.030 161.600 ;
        RECT 18.420 161.400 19.420 161.450 ;
        RECT 20.220 161.200 20.420 162.040 ;
        RECT 20.820 161.600 21.320 161.900 ;
        RECT 21.660 161.600 22.460 161.680 ;
        RECT 20.820 161.450 22.460 161.600 ;
        RECT 20.820 161.400 21.820 161.450 ;
        RECT 22.620 161.200 22.820 162.040 ;
        RECT 23.320 161.600 23.820 161.900 ;
        RECT 24.090 161.600 24.890 161.680 ;
        RECT 23.320 161.450 24.890 161.600 ;
        RECT 23.320 161.400 24.320 161.450 ;
        RECT 25.120 161.200 25.320 162.040 ;
        RECT 25.720 161.600 26.220 161.900 ;
        RECT 26.520 161.600 27.320 161.680 ;
        RECT 25.720 161.450 27.320 161.600 ;
        RECT 25.720 161.400 26.820 161.450 ;
        RECT 27.520 161.200 27.720 162.040 ;
        RECT 28.020 161.900 28.220 163.700 ;
        RECT 30.880 163.400 34.920 163.430 ;
        RECT 38.120 163.400 38.620 163.700 ;
        RECT 30.880 163.200 38.620 163.400 ;
        RECT 28.640 162.400 28.870 163.040 ;
        RECT 28.620 162.040 28.870 162.400 ;
        RECT 36.930 162.300 37.160 163.040 ;
        RECT 37.420 162.300 37.920 162.500 ;
        RECT 36.930 162.040 37.920 162.300 ;
        RECT 28.620 161.900 28.820 162.040 ;
        RECT 28.020 161.600 28.820 161.900 ;
        RECT 37.020 162.000 37.920 162.040 ;
        RECT 30.525 161.600 35.275 161.680 ;
        RECT 28.020 161.450 35.275 161.600 ;
        RECT 28.020 161.400 30.820 161.450 ;
        RECT 37.020 161.200 37.220 162.000 ;
        RECT 8.120 161.000 37.220 161.200 ;
        RECT 2.300 156.310 36.800 156.400 ;
        RECT 2.300 156.200 39.265 156.310 ;
        RECT 2.300 155.700 3.000 156.200 ;
        RECT 6.220 152.665 6.420 156.200 ;
        RECT 6.720 154.140 6.920 156.200 ;
        RECT 7.220 154.575 7.720 155.300 ;
        RECT 7.220 154.400 7.770 154.575 ;
        RECT 7.230 154.345 7.770 154.400 ;
        RECT 6.720 153.800 6.970 154.140 ;
        RECT 6.170 152.400 6.420 152.665 ;
        RECT 6.170 147.975 6.400 152.400 ;
        RECT 6.740 146.140 6.970 153.800 ;
        RECT 8.030 146.400 8.260 154.140 ;
        RECT 8.620 152.665 8.820 156.200 ;
        RECT 12.120 155.500 12.620 156.000 ;
        RECT 9.720 154.575 10.220 155.300 ;
        RECT 9.660 154.400 10.220 154.575 ;
        RECT 12.120 154.600 12.320 155.500 ;
        RECT 12.120 154.530 12.820 154.600 ;
        RECT 12.120 154.400 13.170 154.530 ;
        RECT 9.660 154.345 10.200 154.400 ;
        RECT 12.120 154.140 12.320 154.400 ;
        RECT 12.630 154.300 13.170 154.400 ;
        RECT 8.600 147.975 8.830 152.665 ;
        RECT 9.170 146.400 9.400 154.140 ;
        RECT 8.030 146.200 9.400 146.400 ;
        RECT 8.030 146.140 8.260 146.200 ;
        RECT 9.170 146.140 9.400 146.200 ;
        RECT 10.460 146.400 10.690 154.140 ;
        RECT 12.120 153.900 12.370 154.140 ;
        RECT 11.570 152.600 11.800 152.630 ;
        RECT 11.570 152.400 11.820 152.600 ;
        RECT 11.570 147.960 11.800 152.400 ;
        RECT 12.140 146.400 12.370 153.900 ;
        RECT 10.460 146.200 12.370 146.400 ;
        RECT 10.460 146.140 10.690 146.200 ;
        RECT 12.140 146.140 12.370 146.200 ;
        RECT 13.430 146.400 13.660 154.140 ;
        RECT 14.520 152.665 14.720 156.200 ;
        RECT 15.120 154.140 15.320 156.200 ;
        RECT 15.620 154.575 16.120 155.300 ;
        RECT 15.620 154.400 16.170 154.575 ;
        RECT 15.630 154.345 16.170 154.400 ;
        RECT 15.120 153.800 15.370 154.140 ;
        RECT 14.520 152.400 14.800 152.665 ;
        RECT 14.570 147.975 14.800 152.400 ;
        RECT 13.430 146.140 13.720 146.400 ;
        RECT 15.140 146.140 15.370 153.800 ;
        RECT 16.430 146.400 16.660 154.140 ;
        RECT 17.020 152.670 17.220 156.200 ;
        RECT 20.820 155.500 21.320 156.000 ;
        RECT 18.020 154.600 18.520 155.300 ;
        RECT 18.020 154.400 20.720 154.600 ;
        RECT 21.020 154.545 21.320 155.500 ;
        RECT 21.020 154.400 21.580 154.545 ;
        RECT 18.060 154.350 18.600 154.400 ;
        RECT 20.520 154.155 20.720 154.400 ;
        RECT 21.040 154.315 21.580 154.400 ;
        RECT 17.000 147.980 17.230 152.670 ;
        RECT 17.570 146.400 17.800 154.145 ;
        RECT 16.430 146.200 17.800 146.400 ;
        RECT 16.430 146.140 16.660 146.200 ;
        RECT 17.570 146.145 17.800 146.200 ;
        RECT 18.860 146.400 19.090 154.145 ;
        RECT 20.520 153.900 20.780 154.155 ;
        RECT 19.980 147.975 20.210 152.645 ;
        RECT 20.550 146.400 20.780 153.900 ;
        RECT 18.860 146.200 20.780 146.400 ;
        RECT 18.860 146.145 19.090 146.200 ;
        RECT 20.550 146.155 20.780 146.200 ;
        RECT 21.840 146.400 22.070 154.155 ;
        RECT 22.920 152.665 23.120 156.200 ;
        RECT 23.520 154.140 23.720 156.200 ;
        RECT 24.020 154.575 24.520 155.300 ;
        RECT 24.020 154.400 24.570 154.575 ;
        RECT 24.030 154.345 24.570 154.400 ;
        RECT 23.520 153.800 23.770 154.140 ;
        RECT 22.920 152.400 23.200 152.665 ;
        RECT 22.970 147.975 23.200 152.400 ;
        RECT 21.840 146.155 22.120 146.400 ;
        RECT 13.520 146.100 13.720 146.140 ;
        RECT 13.520 145.900 14.520 146.100 ;
        RECT 13.620 145.400 14.120 145.700 ;
        RECT 14.320 145.600 14.520 145.900 ;
        RECT 14.320 145.400 16.620 145.600 ;
        RECT 6.620 145.200 14.120 145.400 ;
        RECT 6.620 144.040 6.820 145.200 ;
        RECT 7.220 144.430 7.720 145.000 ;
        RECT 7.210 144.200 7.750 144.430 ;
        RECT 9.120 144.040 9.320 145.200 ;
        RECT 9.620 144.430 10.120 145.000 ;
        RECT 9.620 144.300 10.180 144.430 ;
        RECT 9.640 144.200 10.180 144.300 ;
        RECT 11.520 144.040 11.720 145.200 ;
        RECT 12.020 144.430 12.520 145.000 ;
        RECT 12.020 144.300 12.610 144.430 ;
        RECT 12.070 144.200 12.610 144.300 ;
        RECT 13.920 144.040 14.120 145.200 ;
        RECT 16.420 145.000 16.620 145.400 ;
        RECT 18.520 145.400 19.020 145.700 ;
        RECT 21.920 145.400 22.120 146.155 ;
        RECT 23.540 146.140 23.770 153.800 ;
        RECT 24.830 146.500 25.060 154.140 ;
        RECT 25.320 152.665 25.520 156.200 ;
        RECT 26.420 154.575 26.920 155.300 ;
        RECT 26.420 154.400 26.970 154.575 ;
        RECT 26.430 154.345 26.970 154.400 ;
        RECT 25.320 152.400 25.600 152.665 ;
        RECT 25.370 147.975 25.600 152.400 ;
        RECT 25.940 146.500 26.170 154.140 ;
        RECT 24.830 146.300 26.170 146.500 ;
        RECT 24.830 146.140 25.060 146.300 ;
        RECT 25.940 146.140 26.170 146.300 ;
        RECT 27.230 146.400 27.460 154.140 ;
        RECT 27.720 152.665 27.920 156.200 ;
        RECT 28.320 154.140 28.520 156.200 ;
        RECT 28.820 154.575 29.320 155.300 ;
        RECT 28.820 154.400 29.370 154.575 ;
        RECT 28.830 154.345 29.370 154.400 ;
        RECT 28.320 153.800 28.570 154.140 ;
        RECT 27.720 152.400 28.000 152.665 ;
        RECT 27.770 147.975 28.000 152.400 ;
        RECT 27.230 146.140 27.520 146.400 ;
        RECT 28.340 146.140 28.570 153.800 ;
        RECT 29.630 146.400 29.860 154.140 ;
        RECT 30.120 152.665 30.320 156.200 ;
        RECT 31.920 155.500 32.420 156.000 ;
        RECT 31.220 154.575 31.720 155.300 ;
        RECT 31.220 154.400 31.765 154.575 ;
        RECT 31.225 154.345 31.765 154.400 ;
        RECT 32.120 154.140 32.320 155.500 ;
        RECT 30.120 152.400 30.395 152.665 ;
        RECT 30.165 147.975 30.395 152.400 ;
        RECT 30.735 146.400 30.965 154.140 ;
        RECT 29.630 146.200 30.965 146.400 ;
        RECT 29.630 146.140 29.860 146.200 ;
        RECT 30.735 146.140 30.965 146.200 ;
        RECT 32.025 153.900 32.320 154.140 ;
        RECT 32.025 146.140 32.255 153.900 ;
        RECT 32.620 149.980 32.820 156.200 ;
        RECT 36.575 156.080 39.265 156.200 ;
        RECT 33.400 155.800 33.900 156.000 ;
        RECT 33.400 155.740 36.000 155.800 ;
        RECT 33.400 155.600 39.740 155.740 ;
        RECT 33.400 155.500 33.900 155.600 ;
        RECT 35.740 155.510 39.740 155.600 ;
        RECT 39.945 155.300 40.175 155.460 ;
        RECT 40.900 155.300 41.600 155.800 ;
        RECT 33.420 154.800 33.920 155.300 ;
        RECT 39.945 155.100 41.600 155.300 ;
        RECT 41.900 155.100 42.600 155.800 ;
        RECT 39.945 155.000 40.175 155.100 ;
        RECT 33.170 151.700 33.400 152.245 ;
        RECT 33.120 151.365 33.400 151.700 ;
        RECT 33.720 151.860 33.920 154.800 ;
        RECT 35.740 154.800 39.740 154.950 ;
        RECT 43.900 154.800 44.100 180.600 ;
        RECT 60.975 168.500 65.665 168.550 ;
        RECT 71.000 168.500 73.000 210.000 ;
        RECT 48.400 168.000 48.900 168.500 ;
        RECT 60.975 168.320 73.000 168.500 ;
        RECT 65.400 168.300 73.000 168.320 ;
        RECT 56.800 168.000 58.400 168.100 ;
        RECT 69.200 168.000 69.400 168.300 ;
        RECT 48.400 167.640 48.600 168.000 ;
        RECT 49.040 167.900 58.400 168.000 ;
        RECT 66.800 167.980 69.400 168.000 ;
        RECT 49.040 167.770 57.040 167.900 ;
        RECT 48.400 167.500 48.680 167.640 ;
        RECT 48.450 166.840 48.680 167.500 ;
        RECT 57.200 167.500 57.430 167.510 ;
        RECT 57.200 167.000 58.000 167.500 ;
        RECT 57.200 166.970 57.430 167.000 ;
        RECT 49.040 166.600 57.040 166.710 ;
        RECT 35.740 154.720 44.100 154.800 ;
        RECT 39.400 154.600 44.100 154.720 ;
        RECT 38.020 152.500 38.520 153.000 ;
        RECT 38.020 152.250 38.220 152.500 ;
        RECT 35.980 152.020 40.020 152.250 ;
        RECT 33.720 151.600 33.970 151.860 ;
        RECT 42.030 151.700 42.260 151.860 ;
        RECT 33.740 151.440 33.970 151.600 ;
        RECT 42.020 151.440 42.260 151.700 ;
        RECT 33.120 150.900 33.320 151.365 ;
        RECT 42.020 150.900 42.220 151.440 ;
        RECT 33.120 150.700 43.720 150.900 ;
        RECT 39.220 149.995 43.320 150.000 ;
        RECT 32.620 149.500 32.900 149.980 ;
        RECT 35.480 149.800 43.320 149.995 ;
        RECT 35.480 149.765 39.520 149.800 ;
        RECT 33.240 149.500 33.470 149.560 ;
        RECT 32.620 149.300 33.470 149.500 ;
        RECT 41.530 149.400 41.760 149.560 ;
        RECT 32.670 149.080 32.900 149.300 ;
        RECT 33.240 149.140 33.470 149.300 ;
        RECT 41.520 149.200 42.920 149.400 ;
        RECT 41.530 149.140 41.760 149.200 ;
        RECT 42.720 148.000 42.920 149.200 ;
        RECT 42.420 147.700 42.920 148.000 ;
        RECT 41.420 147.640 42.920 147.700 ;
        RECT 33.760 147.500 42.920 147.640 ;
        RECT 33.760 147.410 41.760 147.500 ;
        RECT 33.170 146.800 33.400 147.280 ;
        RECT 41.920 147.100 42.150 147.150 ;
        RECT 43.120 147.100 43.320 149.800 ;
        RECT 41.920 146.900 43.320 147.100 ;
        RECT 33.170 146.480 33.420 146.800 ;
        RECT 41.920 146.610 42.150 146.900 ;
        RECT 42.420 146.600 42.920 146.900 ;
        RECT 27.320 145.400 27.520 146.140 ;
        RECT 33.220 145.800 33.420 146.480 ;
        RECT 33.760 146.120 41.760 146.350 ;
        RECT 33.820 145.800 34.020 146.120 ;
        RECT 43.520 145.800 43.720 150.700 ;
        RECT 33.220 145.600 43.720 145.800 ;
        RECT 18.520 145.200 26.320 145.400 ;
        RECT 27.320 145.200 42.220 145.400 ;
        RECT 14.520 144.430 15.020 145.000 ;
        RECT 16.420 144.800 17.420 145.000 ;
        RECT 14.500 144.200 15.040 144.430 ;
        RECT 16.420 144.040 16.620 144.800 ;
        RECT 16.920 144.430 17.420 144.800 ;
        RECT 16.920 144.300 17.470 144.430 ;
        RECT 16.930 144.200 17.470 144.300 ;
        RECT 18.820 144.040 19.020 145.200 ;
        RECT 19.420 144.430 19.920 145.000 ;
        RECT 19.360 144.300 19.920 144.430 ;
        RECT 19.360 144.200 19.900 144.300 ;
        RECT 21.220 144.040 21.420 145.200 ;
        RECT 21.820 144.430 22.320 145.000 ;
        RECT 21.790 144.200 22.330 144.430 ;
        RECT 23.720 144.040 23.920 145.200 ;
        RECT 24.220 144.430 24.720 145.000 ;
        RECT 24.220 144.200 24.760 144.430 ;
        RECT 26.120 144.040 26.320 145.200 ;
        RECT 26.620 144.430 27.120 145.000 ;
        RECT 26.620 144.300 27.190 144.430 ;
        RECT 26.650 144.200 27.190 144.300 ;
        RECT 32.155 144.300 38.745 144.330 ;
        RECT 42.020 144.300 42.220 145.200 ;
        RECT 32.155 144.100 42.220 144.300 ;
        RECT 6.620 143.800 6.950 144.040 ;
        RECT 6.720 136.040 6.950 143.800 ;
        RECT 8.010 136.300 8.240 144.040 ;
        RECT 9.120 143.800 9.380 144.040 ;
        RECT 8.010 136.040 8.320 136.300 ;
        RECT 9.150 136.040 9.380 143.800 ;
        RECT 10.440 136.300 10.670 144.040 ;
        RECT 11.520 143.800 11.810 144.040 ;
        RECT 10.440 136.040 10.720 136.300 ;
        RECT 11.580 136.040 11.810 143.800 ;
        RECT 12.870 136.300 13.100 144.040 ;
        RECT 13.920 143.800 14.240 144.040 ;
        RECT 12.870 136.040 13.120 136.300 ;
        RECT 14.010 136.040 14.240 143.800 ;
        RECT 15.300 136.300 15.530 144.040 ;
        RECT 16.420 143.800 16.670 144.040 ;
        RECT 15.300 136.040 15.620 136.300 ;
        RECT 16.440 136.040 16.670 143.800 ;
        RECT 17.730 136.300 17.960 144.040 ;
        RECT 18.820 143.800 19.100 144.040 ;
        RECT 17.730 136.040 18.020 136.300 ;
        RECT 18.870 136.040 19.100 143.800 ;
        RECT 20.160 136.300 20.390 144.040 ;
        RECT 21.220 143.800 21.530 144.040 ;
        RECT 20.160 136.040 20.420 136.300 ;
        RECT 21.300 136.040 21.530 143.800 ;
        RECT 22.590 136.040 22.820 144.040 ;
        RECT 23.720 143.800 23.960 144.040 ;
        RECT 23.730 136.040 23.960 143.800 ;
        RECT 25.020 136.300 25.250 144.040 ;
        RECT 26.120 143.800 26.390 144.040 ;
        RECT 25.020 136.040 25.320 136.300 ;
        RECT 26.160 136.040 26.390 143.800 ;
        RECT 27.450 136.300 27.680 144.040 ;
        RECT 42.020 143.940 42.220 144.100 ;
        RECT 28.640 143.200 28.870 143.940 ;
        RECT 42.020 143.600 42.260 143.940 ;
        RECT 28.620 142.940 28.870 143.200 ;
        RECT 42.030 143.200 42.260 143.600 ;
        RECT 42.520 143.200 43.020 143.500 ;
        RECT 42.030 143.000 43.020 143.200 ;
        RECT 42.030 142.940 42.260 143.000 ;
        RECT 28.620 141.640 28.820 142.940 ;
        RECT 31.800 142.350 39.100 142.580 ;
        RECT 30.880 142.000 34.920 142.030 ;
        RECT 38.120 142.000 38.620 142.200 ;
        RECT 30.880 141.800 38.620 142.000 ;
        RECT 38.120 141.700 38.620 141.800 ;
        RECT 38.820 141.800 39.020 142.350 ;
        RECT 43.220 141.800 43.420 145.600 ;
        RECT 28.620 141.300 28.870 141.640 ;
        RECT 28.640 140.640 28.870 141.300 ;
        RECT 36.930 141.000 37.160 141.640 ;
        RECT 38.820 141.600 43.420 141.800 ;
        RECT 37.420 141.000 37.920 141.200 ;
        RECT 36.930 140.700 37.920 141.000 ;
        RECT 36.930 140.640 37.160 140.700 ;
        RECT 38.820 140.500 39.020 141.600 ;
        RECT 37.420 140.300 39.020 140.500 ;
        RECT 35.020 140.280 37.620 140.300 ;
        RECT 30.525 140.200 37.620 140.280 ;
        RECT 28.020 140.100 37.620 140.200 ;
        RECT 28.020 140.050 35.275 140.100 ;
        RECT 28.020 140.000 30.820 140.050 ;
        RECT 28.020 137.900 28.220 140.000 ;
        RECT 30.880 139.700 34.920 139.730 ;
        RECT 38.120 139.700 38.620 140.000 ;
        RECT 30.880 139.500 38.620 139.700 ;
        RECT 28.640 138.700 28.870 139.340 ;
        RECT 28.620 138.340 28.870 138.700 ;
        RECT 36.930 138.700 37.160 139.340 ;
        RECT 37.420 138.700 37.920 138.900 ;
        RECT 36.930 138.400 37.920 138.700 ;
        RECT 36.930 138.340 37.160 138.400 ;
        RECT 28.620 137.900 28.820 138.340 ;
        RECT 30.525 137.900 35.275 137.980 ;
        RECT 28.020 137.750 35.275 137.900 ;
        RECT 28.020 137.700 30.820 137.750 ;
        RECT 27.450 136.040 27.720 136.300 ;
        RECT 6.220 135.600 6.720 135.900 ;
        RECT 7.080 135.600 7.880 135.680 ;
        RECT 6.220 135.450 7.880 135.600 ;
        RECT 6.220 135.400 7.220 135.450 ;
        RECT 8.120 135.200 8.320 136.040 ;
        RECT 8.720 135.600 9.220 135.900 ;
        RECT 9.510 135.600 10.310 135.680 ;
        RECT 8.720 135.450 10.310 135.600 ;
        RECT 8.720 135.400 9.720 135.450 ;
        RECT 10.520 135.200 10.720 136.040 ;
        RECT 11.120 135.600 11.620 135.900 ;
        RECT 11.940 135.600 12.740 135.680 ;
        RECT 11.120 135.450 12.740 135.600 ;
        RECT 11.120 135.400 12.120 135.450 ;
        RECT 12.920 135.200 13.120 136.040 ;
        RECT 13.520 135.600 14.020 135.900 ;
        RECT 14.370 135.600 15.170 135.680 ;
        RECT 13.520 135.450 15.170 135.600 ;
        RECT 13.520 135.400 14.620 135.450 ;
        RECT 15.420 135.200 15.620 136.040 ;
        RECT 15.920 135.600 16.420 135.900 ;
        RECT 16.800 135.600 17.600 135.680 ;
        RECT 17.820 135.600 18.020 136.040 ;
        RECT 15.920 135.400 18.020 135.600 ;
        RECT 18.420 135.600 18.920 135.900 ;
        RECT 19.230 135.600 20.030 135.680 ;
        RECT 18.420 135.450 20.030 135.600 ;
        RECT 18.420 135.400 19.420 135.450 ;
        RECT 20.220 135.200 20.420 136.040 ;
        RECT 20.820 135.600 21.320 135.900 ;
        RECT 21.660 135.600 22.460 135.680 ;
        RECT 20.820 135.450 22.460 135.600 ;
        RECT 20.820 135.400 21.820 135.450 ;
        RECT 22.620 135.200 22.820 136.040 ;
        RECT 23.320 135.600 23.820 135.900 ;
        RECT 24.090 135.600 24.890 135.680 ;
        RECT 23.320 135.450 24.890 135.600 ;
        RECT 23.320 135.400 24.320 135.450 ;
        RECT 25.120 135.200 25.320 136.040 ;
        RECT 25.720 135.600 26.220 135.900 ;
        RECT 26.520 135.600 27.320 135.680 ;
        RECT 25.720 135.450 27.320 135.600 ;
        RECT 25.720 135.400 26.820 135.450 ;
        RECT 27.520 135.200 27.720 136.040 ;
        RECT 28.020 135.900 28.220 137.700 ;
        RECT 30.880 137.400 34.920 137.430 ;
        RECT 38.120 137.400 38.620 137.700 ;
        RECT 30.880 137.200 38.620 137.400 ;
        RECT 28.640 136.400 28.870 137.040 ;
        RECT 28.620 136.040 28.870 136.400 ;
        RECT 36.930 136.300 37.160 137.040 ;
        RECT 37.420 136.300 37.920 136.500 ;
        RECT 36.930 136.040 37.920 136.300 ;
        RECT 28.620 135.900 28.820 136.040 ;
        RECT 28.020 135.600 28.820 135.900 ;
        RECT 37.020 136.000 37.920 136.040 ;
        RECT 30.525 135.600 35.275 135.680 ;
        RECT 28.020 135.450 35.275 135.600 ;
        RECT 28.020 135.400 30.820 135.450 ;
        RECT 37.020 135.200 37.220 136.000 ;
        RECT 8.120 135.000 37.220 135.200 ;
        RECT 43.900 130.800 44.100 154.600 ;
        RECT 48.000 166.480 57.040 166.600 ;
        RECT 48.000 166.400 49.300 166.480 ;
        RECT 48.000 164.200 48.200 166.400 ;
        RECT 48.400 165.500 48.900 166.000 ;
        RECT 58.200 165.600 58.400 167.900 ;
        RECT 59.140 167.800 69.400 167.980 ;
        RECT 59.140 167.750 67.140 167.800 ;
        RECT 67.400 167.490 68.300 167.500 ;
        RECT 67.345 167.000 68.300 167.490 ;
        RECT 67.345 166.950 67.575 167.000 ;
        RECT 59.140 166.460 67.140 166.690 ;
        RECT 56.800 165.570 58.400 165.600 ;
        RECT 48.400 165.210 48.600 165.500 ;
        RECT 49.040 165.400 58.400 165.570 ;
        RECT 59.200 165.550 59.400 166.460 ;
        RECT 60.975 166.100 65.665 166.120 ;
        RECT 69.200 166.100 69.400 167.800 ;
        RECT 60.975 165.900 69.400 166.100 ;
        RECT 60.975 165.890 65.665 165.900 ;
        RECT 49.040 165.340 57.040 165.400 ;
        RECT 48.400 165.000 48.680 165.210 ;
        RECT 57.300 165.080 58.000 165.100 ;
        RECT 48.450 164.410 48.680 165.000 ;
        RECT 57.200 164.600 58.000 165.080 ;
        RECT 57.200 164.540 57.430 164.600 ;
        RECT 49.040 164.200 57.040 164.280 ;
        RECT 48.000 164.050 57.040 164.200 ;
        RECT 48.000 164.000 49.300 164.050 ;
        RECT 48.000 161.800 48.200 164.000 ;
        RECT 48.400 163.100 48.900 163.600 ;
        RECT 58.200 163.200 58.400 165.400 ;
        RECT 59.140 165.320 67.140 165.550 ;
        RECT 67.345 165.000 67.575 165.060 ;
        RECT 67.345 164.520 68.300 165.000 ;
        RECT 67.400 164.500 68.300 164.520 ;
        RECT 59.140 164.030 67.140 164.260 ;
        RECT 56.800 163.140 58.400 163.200 ;
        RECT 48.400 162.780 48.600 163.100 ;
        RECT 49.040 163.000 58.400 163.140 ;
        RECT 49.040 162.910 57.040 163.000 ;
        RECT 48.400 162.600 48.680 162.780 ;
        RECT 57.300 162.650 58.000 162.700 ;
        RECT 48.450 161.980 48.680 162.600 ;
        RECT 57.200 162.200 58.000 162.650 ;
        RECT 57.200 162.110 57.430 162.200 ;
        RECT 49.040 161.800 57.040 161.850 ;
        RECT 48.000 161.620 57.040 161.800 ;
        RECT 48.000 161.600 49.300 161.620 ;
        RECT 48.000 159.300 48.200 161.600 ;
        RECT 48.400 160.700 48.900 161.200 ;
        RECT 58.200 161.100 58.400 163.000 ;
        RECT 59.200 162.580 59.400 164.030 ;
        RECT 60.960 162.920 65.630 163.150 ;
        RECT 65.400 162.900 65.600 162.920 ;
        RECT 66.900 162.580 69.000 162.600 ;
        RECT 59.140 162.400 69.000 162.580 ;
        RECT 59.140 162.350 67.140 162.400 ;
        RECT 67.400 162.090 67.600 162.400 ;
        RECT 68.500 162.100 69.000 162.400 ;
        RECT 67.300 161.900 67.600 162.090 ;
        RECT 67.300 161.550 67.530 161.900 ;
        RECT 59.140 161.200 67.140 161.290 ;
        RECT 58.200 160.800 58.700 161.100 ;
        RECT 56.800 160.710 58.700 160.800 ;
        RECT 48.400 160.350 48.600 160.700 ;
        RECT 49.040 160.600 58.700 160.710 ;
        RECT 58.900 161.060 67.140 161.200 ;
        RECT 58.900 161.000 59.400 161.060 ;
        RECT 49.040 160.480 57.040 160.600 ;
        RECT 58.900 160.400 59.100 161.000 ;
        RECT 48.400 160.100 48.680 160.350 ;
        RECT 48.450 159.550 48.680 160.100 ;
        RECT 57.200 160.200 57.430 160.220 ;
        RECT 58.400 160.200 59.100 160.400 ;
        RECT 69.200 160.200 69.400 165.900 ;
        RECT 57.200 159.700 58.000 160.200 ;
        RECT 57.200 159.680 57.430 159.700 ;
        RECT 49.040 159.300 57.040 159.420 ;
        RECT 48.000 159.190 57.040 159.300 ;
        RECT 48.000 159.100 49.300 159.190 ;
        RECT 48.000 154.500 48.200 159.100 ;
        RECT 48.400 158.300 48.900 158.800 ;
        RECT 58.400 158.300 58.600 160.200 ;
        RECT 65.400 160.150 69.400 160.200 ;
        RECT 60.975 160.000 69.400 160.150 ;
        RECT 60.975 159.920 65.665 160.000 ;
        RECT 69.200 159.600 69.400 160.000 ;
        RECT 66.800 159.580 69.400 159.600 ;
        RECT 59.140 159.400 69.400 159.580 ;
        RECT 59.140 159.350 67.140 159.400 ;
        RECT 67.400 159.090 68.300 159.100 ;
        RECT 67.345 158.600 68.300 159.090 ;
        RECT 67.345 158.550 67.575 158.600 ;
        RECT 48.400 157.920 48.600 158.300 ;
        RECT 56.800 158.280 58.600 158.300 ;
        RECT 49.040 158.100 58.600 158.280 ;
        RECT 49.040 158.050 57.040 158.100 ;
        RECT 48.400 157.120 48.680 157.920 ;
        RECT 57.800 157.800 58.000 158.100 ;
        RECT 59.140 158.060 67.140 158.290 ;
        RECT 57.300 157.790 58.000 157.800 ;
        RECT 57.200 157.300 58.000 157.790 ;
        RECT 57.200 157.250 57.430 157.300 ;
        RECT 59.200 157.150 59.400 158.060 ;
        RECT 60.980 157.700 65.670 157.720 ;
        RECT 69.200 157.700 69.400 159.400 ;
        RECT 60.980 157.500 69.400 157.700 ;
        RECT 60.980 157.490 65.670 157.500 ;
        RECT 48.400 156.900 48.600 157.120 ;
        RECT 49.040 156.900 57.040 156.990 ;
        RECT 59.145 156.920 67.145 157.150 ;
        RECT 48.400 156.760 57.040 156.900 ;
        RECT 48.400 156.700 49.300 156.760 ;
        RECT 67.400 156.660 68.300 156.700 ;
        RECT 48.400 155.800 48.900 156.300 ;
        RECT 67.350 156.200 68.300 156.660 ;
        RECT 58.200 155.900 58.700 156.200 ;
        RECT 67.350 156.120 67.600 156.200 ;
        RECT 56.800 155.850 58.700 155.900 ;
        RECT 48.400 155.490 48.600 155.800 ;
        RECT 49.040 155.700 58.700 155.850 ;
        RECT 49.040 155.620 57.040 155.700 ;
        RECT 48.400 155.300 48.680 155.490 ;
        RECT 48.450 154.690 48.680 155.300 ;
        RECT 57.200 155.300 57.430 155.360 ;
        RECT 57.200 154.820 58.000 155.300 ;
        RECT 57.300 154.800 58.000 154.820 ;
        RECT 49.040 154.500 57.040 154.560 ;
        RECT 48.000 154.330 57.040 154.500 ;
        RECT 48.000 154.300 49.300 154.330 ;
        RECT 48.000 152.100 48.200 154.300 ;
        RECT 48.400 153.400 48.900 153.900 ;
        RECT 58.200 153.500 58.400 155.700 ;
        RECT 59.145 155.630 67.145 155.860 ;
        RECT 59.200 154.170 59.400 155.630 ;
        RECT 60.975 154.510 65.645 154.740 ;
        RECT 67.400 154.200 67.600 156.120 ;
        RECT 66.900 154.170 67.600 154.200 ;
        RECT 59.155 154.000 67.600 154.170 ;
        RECT 59.155 153.940 67.155 154.000 ;
        RECT 68.500 153.700 69.000 153.900 ;
        RECT 67.400 153.680 69.000 153.700 ;
        RECT 56.800 153.420 58.400 153.500 ;
        RECT 48.400 153.060 48.600 153.400 ;
        RECT 49.040 153.300 58.400 153.420 ;
        RECT 49.040 153.190 57.040 153.300 ;
        RECT 48.400 152.900 48.680 153.060 ;
        RECT 48.450 152.260 48.680 152.900 ;
        RECT 57.200 152.900 57.430 152.930 ;
        RECT 57.200 152.400 58.000 152.900 ;
        RECT 58.200 152.800 58.400 153.300 ;
        RECT 67.315 153.400 69.000 153.680 ;
        RECT 67.315 153.140 67.545 153.400 ;
        RECT 59.155 152.800 67.155 152.880 ;
        RECT 58.200 152.650 67.155 152.800 ;
        RECT 58.200 152.600 59.400 152.650 ;
        RECT 57.200 152.390 57.430 152.400 ;
        RECT 49.040 152.100 57.040 152.130 ;
        RECT 48.000 151.900 57.040 152.100 ;
        RECT 48.000 149.600 48.200 151.900 ;
        RECT 48.400 150.900 48.900 151.400 ;
        RECT 58.200 151.000 58.400 152.600 ;
        RECT 69.200 151.800 69.400 157.500 ;
        RECT 65.400 151.750 69.400 151.800 ;
        RECT 60.975 151.600 69.400 151.750 ;
        RECT 60.975 151.520 65.665 151.600 ;
        RECT 69.200 151.200 69.400 151.600 ;
        RECT 66.800 151.180 69.400 151.200 ;
        RECT 56.800 150.990 58.400 151.000 ;
        RECT 48.400 150.630 48.600 150.900 ;
        RECT 49.040 150.800 58.400 150.990 ;
        RECT 59.140 151.000 69.400 151.180 ;
        RECT 59.140 150.950 67.140 151.000 ;
        RECT 49.040 150.760 57.040 150.800 ;
        RECT 48.400 150.400 48.680 150.630 ;
        RECT 48.450 149.830 48.680 150.400 ;
        RECT 57.200 150.000 58.000 150.500 ;
        RECT 57.200 149.960 57.430 150.000 ;
        RECT 49.040 149.600 57.040 149.700 ;
        RECT 48.000 149.470 57.040 149.600 ;
        RECT 48.000 149.400 49.300 149.470 ;
        RECT 48.000 147.200 48.200 149.400 ;
        RECT 48.400 148.500 48.900 149.000 ;
        RECT 58.200 148.600 58.400 150.800 ;
        RECT 67.400 150.690 68.300 150.700 ;
        RECT 67.345 150.200 68.300 150.690 ;
        RECT 67.345 150.150 67.575 150.200 ;
        RECT 59.140 149.660 67.140 149.890 ;
        RECT 59.300 148.780 59.500 149.660 ;
        RECT 69.200 149.400 69.400 151.000 ;
        RECT 65.400 149.350 69.400 149.400 ;
        RECT 60.975 149.200 69.400 149.350 ;
        RECT 60.975 149.120 65.665 149.200 ;
        RECT 56.800 148.560 58.400 148.600 ;
        RECT 48.400 148.200 48.600 148.500 ;
        RECT 49.040 148.400 58.400 148.560 ;
        RECT 59.140 148.550 67.140 148.780 ;
        RECT 49.040 148.330 57.040 148.400 ;
        RECT 67.400 148.290 68.300 148.300 ;
        RECT 48.400 147.900 48.680 148.200 ;
        RECT 57.300 148.070 58.000 148.100 ;
        RECT 48.450 147.400 48.680 147.900 ;
        RECT 57.200 147.600 58.000 148.070 ;
        RECT 67.345 147.800 68.300 148.290 ;
        RECT 67.345 147.750 67.575 147.800 ;
        RECT 57.200 147.530 57.430 147.600 ;
        RECT 59.140 147.400 67.140 147.490 ;
        RECT 49.040 147.200 57.040 147.270 ;
        RECT 48.000 147.040 57.040 147.200 ;
        RECT 58.200 147.260 67.140 147.400 ;
        RECT 58.200 147.200 59.400 147.260 ;
        RECT 48.000 147.000 49.300 147.040 ;
        RECT 48.000 137.700 48.200 147.000 ;
        RECT 48.400 146.500 53.200 146.700 ;
        RECT 48.400 146.100 48.900 146.500 ;
        RECT 50.700 146.100 50.900 146.500 ;
        RECT 48.400 146.080 49.400 146.100 ;
        RECT 50.700 146.080 51.700 146.100 ;
        RECT 48.400 145.900 50.040 146.080 ;
        RECT 48.400 144.195 48.600 145.900 ;
        RECT 49.040 145.850 50.040 145.900 ;
        RECT 50.700 145.900 52.340 146.080 ;
        RECT 50.700 144.195 50.900 145.900 ;
        RECT 51.340 145.850 52.340 145.900 ;
        RECT 53.000 144.195 53.200 146.500 ;
        RECT 54.300 146.080 56.200 146.100 ;
        RECT 53.640 145.900 56.940 146.080 ;
        RECT 53.640 145.850 54.640 145.900 ;
        RECT 55.940 145.850 56.940 145.900 ;
        RECT 48.400 143.900 48.680 144.195 ;
        RECT 50.700 143.900 50.980 144.195 ;
        RECT 53.000 143.900 53.280 144.195 ;
        RECT 48.450 139.445 48.680 143.900 ;
        RECT 50.200 139.800 50.430 143.840 ;
        RECT 49.040 137.700 50.040 137.790 ;
        RECT 48.000 137.560 50.040 137.700 ;
        RECT 48.000 137.500 49.300 137.560 ;
        RECT 49.000 137.300 49.300 137.500 ;
        RECT 49.000 136.800 49.500 137.300 ;
        RECT 50.200 136.600 50.400 139.800 ;
        RECT 50.750 139.445 50.980 143.900 ;
        RECT 52.500 139.800 52.730 143.840 ;
        RECT 51.340 137.560 52.340 137.790 ;
        RECT 51.400 137.300 51.700 137.560 ;
        RECT 51.400 136.800 51.900 137.300 ;
        RECT 52.500 136.600 52.700 139.800 ;
        RECT 53.050 139.700 53.280 143.900 ;
        RECT 54.800 139.800 55.030 143.840 ;
        RECT 53.050 139.445 53.300 139.700 ;
        RECT 53.100 137.300 53.300 139.445 ;
        RECT 53.640 137.560 54.640 137.790 ;
        RECT 53.700 137.300 54.000 137.560 ;
        RECT 53.100 137.100 53.500 137.300 ;
        RECT 50.200 136.100 50.700 136.600 ;
        RECT 52.500 136.100 53.000 136.600 ;
        RECT 53.300 135.900 53.500 137.100 ;
        RECT 53.700 136.800 54.200 137.300 ;
        RECT 54.800 136.600 55.000 139.800 ;
        RECT 54.700 136.100 55.200 136.600 ;
        RECT 55.350 135.900 55.580 142.920 ;
        RECT 53.300 135.700 55.580 135.900 ;
        RECT 54.600 131.500 54.800 135.700 ;
        RECT 55.350 135.620 55.580 135.700 ;
        RECT 57.100 135.975 57.330 142.565 ;
        RECT 57.100 132.700 57.300 135.975 ;
        RECT 58.200 132.700 58.400 147.200 ;
        RECT 69.200 147.000 69.400 149.200 ;
        RECT 65.400 146.950 69.400 147.000 ;
        RECT 60.975 146.800 69.400 146.950 ;
        RECT 60.975 146.720 65.665 146.800 ;
        RECT 69.200 146.400 69.400 146.800 ;
        RECT 66.800 146.380 69.400 146.400 ;
        RECT 59.140 146.200 69.400 146.380 ;
        RECT 59.140 146.150 67.140 146.200 ;
        RECT 67.400 145.890 68.300 145.900 ;
        RECT 67.345 145.400 68.300 145.890 ;
        RECT 67.345 145.350 67.575 145.400 ;
        RECT 59.140 144.860 67.140 145.090 ;
        RECT 59.200 143.985 59.400 144.860 ;
        RECT 69.200 144.600 69.400 146.200 ;
        RECT 65.400 144.555 69.400 144.600 ;
        RECT 60.975 144.400 69.400 144.555 ;
        RECT 60.975 144.325 65.665 144.400 ;
        RECT 59.140 143.755 67.140 143.985 ;
        RECT 67.400 143.495 68.300 143.500 ;
        RECT 67.345 143.000 68.300 143.495 ;
        RECT 67.345 142.955 67.575 143.000 ;
        RECT 59.140 142.600 67.140 142.695 ;
        RECT 68.500 142.600 69.000 142.800 ;
        RECT 59.140 142.465 69.000 142.600 ;
        RECT 66.900 142.400 69.000 142.465 ;
        RECT 68.500 142.300 69.000 142.400 ;
        RECT 69.200 142.100 69.400 144.400 ;
        RECT 62.300 142.050 69.400 142.100 ;
        RECT 62.080 141.900 69.400 142.050 ;
        RECT 62.080 141.820 62.980 141.900 ;
        RECT 59.480 141.500 60.280 141.550 ;
        RECT 56.600 132.690 58.400 132.700 ;
        RECT 55.940 132.500 58.400 132.690 ;
        RECT 58.600 141.320 60.280 141.500 ;
        RECT 62.300 141.480 62.500 141.820 ;
        RECT 63.700 141.550 64.700 141.600 ;
        RECT 58.600 141.300 59.800 141.320 ;
        RECT 58.600 140.900 58.800 141.300 ;
        RECT 62.140 141.250 62.560 141.480 ;
        RECT 63.700 141.400 65.245 141.550 ;
        RECT 59.120 140.900 59.350 140.960 ;
        RECT 58.600 140.700 59.350 140.900 ;
        RECT 55.940 132.460 56.940 132.500 ;
        RECT 56.000 132.200 56.200 132.460 ;
        RECT 56.000 131.700 56.500 132.200 ;
        RECT 58.600 131.500 58.800 140.700 ;
        RECT 59.120 132.960 59.350 140.700 ;
        RECT 60.410 133.300 60.640 140.960 ;
        RECT 62.765 135.500 62.995 139.240 ;
        RECT 62.765 135.200 63.000 135.500 ;
        RECT 60.410 132.960 60.700 133.300 ;
        RECT 62.200 133.190 62.400 133.200 ;
        RECT 62.140 132.960 62.560 133.190 ;
        RECT 59.610 132.570 60.150 132.800 ;
        RECT 59.900 132.300 60.100 132.570 ;
        RECT 59.600 131.800 60.100 132.300 ;
        RECT 60.500 132.300 60.700 132.960 ;
        RECT 60.500 132.000 61.000 132.300 ;
        RECT 62.200 132.000 62.400 132.960 ;
        RECT 60.500 131.800 62.400 132.000 ;
        RECT 54.600 131.300 58.800 131.500 ;
        RECT 59.900 131.600 60.100 131.800 ;
        RECT 62.800 131.600 63.000 135.200 ;
        RECT 59.900 131.400 63.000 131.600 ;
        RECT 63.700 132.700 63.900 141.400 ;
        RECT 64.365 141.320 65.245 141.400 ;
        RECT 67.800 141.000 68.300 141.300 ;
        RECT 64.600 140.980 68.300 141.000 ;
        RECT 64.440 140.800 68.300 140.980 ;
        RECT 68.500 140.800 69.000 141.300 ;
        RECT 64.440 140.750 64.860 140.800 ;
        RECT 68.600 139.100 68.800 140.800 ;
        RECT 65.020 136.700 65.250 138.740 ;
        RECT 65.020 136.500 66.000 136.700 ;
        RECT 65.020 134.700 65.250 136.500 ;
        RECT 65.500 136.200 66.000 136.500 ;
        RECT 67.720 135.400 67.950 139.100 ;
        RECT 67.600 135.100 67.950 135.400 ;
        RECT 68.510 138.800 68.800 139.100 ;
        RECT 68.510 135.100 68.740 138.800 ;
        RECT 69.200 138.265 69.400 141.900 ;
        RECT 69.080 137.900 69.400 138.265 ;
        RECT 69.080 135.575 69.310 137.900 ;
        RECT 63.700 132.690 64.700 132.700 ;
        RECT 63.700 132.500 64.860 132.690 ;
        RECT 58.600 131.200 58.800 131.300 ;
        RECT 63.700 131.200 63.900 132.500 ;
        RECT 64.440 132.460 64.860 132.500 ;
        RECT 58.600 131.000 63.900 131.200 ;
        RECT 67.600 130.800 67.800 135.100 ;
        RECT 68.000 134.665 68.460 134.895 ;
        RECT 68.100 133.900 68.300 134.665 ;
        RECT 68.100 133.200 68.800 133.900 ;
        RECT 68.100 132.200 68.800 132.900 ;
        RECT 43.900 130.600 67.800 130.800 ;
        RECT 2.300 130.310 36.800 130.400 ;
        RECT 2.300 130.200 39.265 130.310 ;
        RECT 2.300 129.700 3.000 130.200 ;
        RECT 6.220 126.665 6.420 130.200 ;
        RECT 6.720 128.140 6.920 130.200 ;
        RECT 7.220 128.575 7.720 129.300 ;
        RECT 7.220 128.400 7.770 128.575 ;
        RECT 7.230 128.345 7.770 128.400 ;
        RECT 6.720 127.800 6.970 128.140 ;
        RECT 6.170 126.400 6.420 126.665 ;
        RECT 6.170 121.975 6.400 126.400 ;
        RECT 6.740 120.140 6.970 127.800 ;
        RECT 8.030 120.400 8.260 128.140 ;
        RECT 8.620 126.665 8.820 130.200 ;
        RECT 12.120 129.500 12.620 130.000 ;
        RECT 9.720 128.575 10.220 129.300 ;
        RECT 9.660 128.400 10.220 128.575 ;
        RECT 12.120 128.600 12.320 129.500 ;
        RECT 12.120 128.530 12.820 128.600 ;
        RECT 12.120 128.400 13.170 128.530 ;
        RECT 9.660 128.345 10.200 128.400 ;
        RECT 12.120 128.140 12.320 128.400 ;
        RECT 12.630 128.300 13.170 128.400 ;
        RECT 8.600 121.975 8.830 126.665 ;
        RECT 9.170 120.400 9.400 128.140 ;
        RECT 8.030 120.200 9.400 120.400 ;
        RECT 8.030 120.140 8.260 120.200 ;
        RECT 9.170 120.140 9.400 120.200 ;
        RECT 10.460 120.400 10.690 128.140 ;
        RECT 12.120 127.900 12.370 128.140 ;
        RECT 11.570 126.600 11.800 126.630 ;
        RECT 11.570 126.400 11.820 126.600 ;
        RECT 11.570 121.960 11.800 126.400 ;
        RECT 12.140 120.400 12.370 127.900 ;
        RECT 10.460 120.200 12.370 120.400 ;
        RECT 10.460 120.140 10.690 120.200 ;
        RECT 12.140 120.140 12.370 120.200 ;
        RECT 13.430 120.400 13.660 128.140 ;
        RECT 14.520 126.665 14.720 130.200 ;
        RECT 15.120 128.140 15.320 130.200 ;
        RECT 15.620 128.575 16.120 129.300 ;
        RECT 15.620 128.400 16.170 128.575 ;
        RECT 15.630 128.345 16.170 128.400 ;
        RECT 15.120 127.800 15.370 128.140 ;
        RECT 14.520 126.400 14.800 126.665 ;
        RECT 14.570 121.975 14.800 126.400 ;
        RECT 13.430 120.140 13.720 120.400 ;
        RECT 15.140 120.140 15.370 127.800 ;
        RECT 16.430 120.400 16.660 128.140 ;
        RECT 17.020 126.670 17.220 130.200 ;
        RECT 20.820 129.500 21.320 130.000 ;
        RECT 18.020 128.600 18.520 129.300 ;
        RECT 18.020 128.400 20.720 128.600 ;
        RECT 21.020 128.545 21.320 129.500 ;
        RECT 21.020 128.400 21.580 128.545 ;
        RECT 18.060 128.350 18.600 128.400 ;
        RECT 20.520 128.155 20.720 128.400 ;
        RECT 21.040 128.315 21.580 128.400 ;
        RECT 17.000 121.980 17.230 126.670 ;
        RECT 17.570 120.400 17.800 128.145 ;
        RECT 16.430 120.200 17.800 120.400 ;
        RECT 16.430 120.140 16.660 120.200 ;
        RECT 17.570 120.145 17.800 120.200 ;
        RECT 18.860 120.400 19.090 128.145 ;
        RECT 20.520 127.900 20.780 128.155 ;
        RECT 19.980 121.975 20.210 126.645 ;
        RECT 20.550 120.400 20.780 127.900 ;
        RECT 18.860 120.200 20.780 120.400 ;
        RECT 18.860 120.145 19.090 120.200 ;
        RECT 20.550 120.155 20.780 120.200 ;
        RECT 21.840 120.400 22.070 128.155 ;
        RECT 22.920 126.665 23.120 130.200 ;
        RECT 23.520 128.140 23.720 130.200 ;
        RECT 24.020 128.575 24.520 129.300 ;
        RECT 24.020 128.400 24.570 128.575 ;
        RECT 24.030 128.345 24.570 128.400 ;
        RECT 23.520 127.800 23.770 128.140 ;
        RECT 22.920 126.400 23.200 126.665 ;
        RECT 22.970 121.975 23.200 126.400 ;
        RECT 21.840 120.155 22.120 120.400 ;
        RECT 13.520 120.100 13.720 120.140 ;
        RECT 13.520 119.900 14.520 120.100 ;
        RECT 13.620 119.400 14.120 119.700 ;
        RECT 14.320 119.600 14.520 119.900 ;
        RECT 14.320 119.400 16.620 119.600 ;
        RECT 6.620 119.200 14.120 119.400 ;
        RECT 6.620 118.040 6.820 119.200 ;
        RECT 7.220 118.430 7.720 119.000 ;
        RECT 7.210 118.200 7.750 118.430 ;
        RECT 9.120 118.040 9.320 119.200 ;
        RECT 9.620 118.430 10.120 119.000 ;
        RECT 9.620 118.300 10.180 118.430 ;
        RECT 9.640 118.200 10.180 118.300 ;
        RECT 11.520 118.040 11.720 119.200 ;
        RECT 12.020 118.430 12.520 119.000 ;
        RECT 12.020 118.300 12.610 118.430 ;
        RECT 12.070 118.200 12.610 118.300 ;
        RECT 13.920 118.040 14.120 119.200 ;
        RECT 16.420 119.000 16.620 119.400 ;
        RECT 18.520 119.400 19.020 119.700 ;
        RECT 21.920 119.400 22.120 120.155 ;
        RECT 23.540 120.140 23.770 127.800 ;
        RECT 24.830 120.500 25.060 128.140 ;
        RECT 25.320 126.665 25.520 130.200 ;
        RECT 26.420 128.575 26.920 129.300 ;
        RECT 26.420 128.400 26.970 128.575 ;
        RECT 26.430 128.345 26.970 128.400 ;
        RECT 25.320 126.400 25.600 126.665 ;
        RECT 25.370 121.975 25.600 126.400 ;
        RECT 25.940 120.500 26.170 128.140 ;
        RECT 24.830 120.300 26.170 120.500 ;
        RECT 24.830 120.140 25.060 120.300 ;
        RECT 25.940 120.140 26.170 120.300 ;
        RECT 27.230 120.400 27.460 128.140 ;
        RECT 27.720 126.665 27.920 130.200 ;
        RECT 28.320 128.140 28.520 130.200 ;
        RECT 28.820 128.575 29.320 129.300 ;
        RECT 28.820 128.400 29.370 128.575 ;
        RECT 28.830 128.345 29.370 128.400 ;
        RECT 28.320 127.800 28.570 128.140 ;
        RECT 27.720 126.400 28.000 126.665 ;
        RECT 27.770 121.975 28.000 126.400 ;
        RECT 27.230 120.140 27.520 120.400 ;
        RECT 28.340 120.140 28.570 127.800 ;
        RECT 29.630 120.400 29.860 128.140 ;
        RECT 30.120 126.665 30.320 130.200 ;
        RECT 31.920 129.500 32.420 130.000 ;
        RECT 31.220 128.575 31.720 129.300 ;
        RECT 31.220 128.400 31.765 128.575 ;
        RECT 31.225 128.345 31.765 128.400 ;
        RECT 32.120 128.140 32.320 129.500 ;
        RECT 30.120 126.400 30.395 126.665 ;
        RECT 30.165 121.975 30.395 126.400 ;
        RECT 30.735 120.400 30.965 128.140 ;
        RECT 29.630 120.200 30.965 120.400 ;
        RECT 29.630 120.140 29.860 120.200 ;
        RECT 30.735 120.140 30.965 120.200 ;
        RECT 32.025 127.900 32.320 128.140 ;
        RECT 32.025 120.140 32.255 127.900 ;
        RECT 32.620 123.980 32.820 130.200 ;
        RECT 36.575 130.080 39.265 130.200 ;
        RECT 33.400 129.800 33.900 130.000 ;
        RECT 33.400 129.740 36.000 129.800 ;
        RECT 33.400 129.600 39.740 129.740 ;
        RECT 33.400 129.500 33.900 129.600 ;
        RECT 35.740 129.510 39.740 129.600 ;
        RECT 39.945 129.300 40.175 129.460 ;
        RECT 40.900 129.300 41.600 129.800 ;
        RECT 33.420 128.800 33.920 129.300 ;
        RECT 39.945 129.100 41.600 129.300 ;
        RECT 41.900 129.100 42.600 129.800 ;
        RECT 39.945 129.000 40.175 129.100 ;
        RECT 33.170 125.700 33.400 126.245 ;
        RECT 33.120 125.365 33.400 125.700 ;
        RECT 33.720 125.860 33.920 128.800 ;
        RECT 35.740 128.800 39.740 128.950 ;
        RECT 43.900 128.800 44.100 130.600 ;
        RECT 35.740 128.720 44.100 128.800 ;
        RECT 39.400 128.600 44.100 128.720 ;
        RECT 38.020 126.500 38.520 127.000 ;
        RECT 38.020 126.250 38.220 126.500 ;
        RECT 35.980 126.020 40.020 126.250 ;
        RECT 33.720 125.600 33.970 125.860 ;
        RECT 42.030 125.700 42.260 125.860 ;
        RECT 33.740 125.440 33.970 125.600 ;
        RECT 42.020 125.440 42.260 125.700 ;
        RECT 33.120 124.900 33.320 125.365 ;
        RECT 42.020 124.900 42.220 125.440 ;
        RECT 33.120 124.700 43.720 124.900 ;
        RECT 39.220 123.995 43.320 124.000 ;
        RECT 32.620 123.500 32.900 123.980 ;
        RECT 35.480 123.800 43.320 123.995 ;
        RECT 35.480 123.765 39.520 123.800 ;
        RECT 33.240 123.500 33.470 123.560 ;
        RECT 32.620 123.300 33.470 123.500 ;
        RECT 41.530 123.400 41.760 123.560 ;
        RECT 32.670 123.080 32.900 123.300 ;
        RECT 33.240 123.140 33.470 123.300 ;
        RECT 41.520 123.200 42.920 123.400 ;
        RECT 41.530 123.140 41.760 123.200 ;
        RECT 42.720 122.000 42.920 123.200 ;
        RECT 42.420 121.700 42.920 122.000 ;
        RECT 41.420 121.640 42.920 121.700 ;
        RECT 33.760 121.500 42.920 121.640 ;
        RECT 33.760 121.410 41.760 121.500 ;
        RECT 33.170 120.800 33.400 121.280 ;
        RECT 41.920 121.100 42.150 121.150 ;
        RECT 43.120 121.100 43.320 123.800 ;
        RECT 41.920 120.900 43.320 121.100 ;
        RECT 33.170 120.480 33.420 120.800 ;
        RECT 41.920 120.610 42.150 120.900 ;
        RECT 42.420 120.600 42.920 120.900 ;
        RECT 27.320 119.400 27.520 120.140 ;
        RECT 33.220 119.800 33.420 120.480 ;
        RECT 33.760 120.120 41.760 120.350 ;
        RECT 33.820 119.800 34.020 120.120 ;
        RECT 43.520 119.800 43.720 124.700 ;
        RECT 33.220 119.600 43.720 119.800 ;
        RECT 18.520 119.200 26.320 119.400 ;
        RECT 27.320 119.200 42.220 119.400 ;
        RECT 14.520 118.430 15.020 119.000 ;
        RECT 16.420 118.800 17.420 119.000 ;
        RECT 14.500 118.200 15.040 118.430 ;
        RECT 16.420 118.040 16.620 118.800 ;
        RECT 16.920 118.430 17.420 118.800 ;
        RECT 16.920 118.300 17.470 118.430 ;
        RECT 16.930 118.200 17.470 118.300 ;
        RECT 18.820 118.040 19.020 119.200 ;
        RECT 19.420 118.430 19.920 119.000 ;
        RECT 19.360 118.300 19.920 118.430 ;
        RECT 19.360 118.200 19.900 118.300 ;
        RECT 21.220 118.040 21.420 119.200 ;
        RECT 21.820 118.430 22.320 119.000 ;
        RECT 21.790 118.200 22.330 118.430 ;
        RECT 23.720 118.040 23.920 119.200 ;
        RECT 24.220 118.430 24.720 119.000 ;
        RECT 24.220 118.200 24.760 118.430 ;
        RECT 26.120 118.040 26.320 119.200 ;
        RECT 26.620 118.430 27.120 119.000 ;
        RECT 26.620 118.300 27.190 118.430 ;
        RECT 26.650 118.200 27.190 118.300 ;
        RECT 32.155 118.300 38.745 118.330 ;
        RECT 42.020 118.300 42.220 119.200 ;
        RECT 32.155 118.100 42.220 118.300 ;
        RECT 6.620 117.800 6.950 118.040 ;
        RECT 6.720 110.040 6.950 117.800 ;
        RECT 8.010 110.300 8.240 118.040 ;
        RECT 9.120 117.800 9.380 118.040 ;
        RECT 8.010 110.040 8.320 110.300 ;
        RECT 9.150 110.040 9.380 117.800 ;
        RECT 10.440 110.300 10.670 118.040 ;
        RECT 11.520 117.800 11.810 118.040 ;
        RECT 10.440 110.040 10.720 110.300 ;
        RECT 11.580 110.040 11.810 117.800 ;
        RECT 12.870 110.300 13.100 118.040 ;
        RECT 13.920 117.800 14.240 118.040 ;
        RECT 12.870 110.040 13.120 110.300 ;
        RECT 14.010 110.040 14.240 117.800 ;
        RECT 15.300 110.300 15.530 118.040 ;
        RECT 16.420 117.800 16.670 118.040 ;
        RECT 15.300 110.040 15.620 110.300 ;
        RECT 16.440 110.040 16.670 117.800 ;
        RECT 17.730 110.300 17.960 118.040 ;
        RECT 18.820 117.800 19.100 118.040 ;
        RECT 17.730 110.040 18.020 110.300 ;
        RECT 18.870 110.040 19.100 117.800 ;
        RECT 20.160 110.300 20.390 118.040 ;
        RECT 21.220 117.800 21.530 118.040 ;
        RECT 20.160 110.040 20.420 110.300 ;
        RECT 21.300 110.040 21.530 117.800 ;
        RECT 22.590 110.040 22.820 118.040 ;
        RECT 23.720 117.800 23.960 118.040 ;
        RECT 23.730 110.040 23.960 117.800 ;
        RECT 25.020 110.300 25.250 118.040 ;
        RECT 26.120 117.800 26.390 118.040 ;
        RECT 25.020 110.040 25.320 110.300 ;
        RECT 26.160 110.040 26.390 117.800 ;
        RECT 27.450 110.300 27.680 118.040 ;
        RECT 42.020 117.940 42.220 118.100 ;
        RECT 28.640 117.200 28.870 117.940 ;
        RECT 42.020 117.600 42.260 117.940 ;
        RECT 28.620 116.940 28.870 117.200 ;
        RECT 42.030 117.200 42.260 117.600 ;
        RECT 42.520 117.200 43.020 117.500 ;
        RECT 42.030 117.000 43.020 117.200 ;
        RECT 42.030 116.940 42.260 117.000 ;
        RECT 28.620 115.640 28.820 116.940 ;
        RECT 31.800 116.350 39.100 116.580 ;
        RECT 30.880 116.000 34.920 116.030 ;
        RECT 38.120 116.000 38.620 116.200 ;
        RECT 30.880 115.800 38.620 116.000 ;
        RECT 38.120 115.700 38.620 115.800 ;
        RECT 38.820 115.800 39.020 116.350 ;
        RECT 43.220 115.800 43.420 119.600 ;
        RECT 28.620 115.300 28.870 115.640 ;
        RECT 28.640 114.640 28.870 115.300 ;
        RECT 36.930 115.000 37.160 115.640 ;
        RECT 38.820 115.600 43.420 115.800 ;
        RECT 37.420 115.000 37.920 115.200 ;
        RECT 36.930 114.700 37.920 115.000 ;
        RECT 36.930 114.640 37.160 114.700 ;
        RECT 38.820 114.500 39.020 115.600 ;
        RECT 37.420 114.300 39.020 114.500 ;
        RECT 35.020 114.280 37.620 114.300 ;
        RECT 30.525 114.200 37.620 114.280 ;
        RECT 28.020 114.100 37.620 114.200 ;
        RECT 28.020 114.050 35.275 114.100 ;
        RECT 28.020 114.000 30.820 114.050 ;
        RECT 28.020 111.900 28.220 114.000 ;
        RECT 30.880 113.700 34.920 113.730 ;
        RECT 38.120 113.700 38.620 114.000 ;
        RECT 30.880 113.500 38.620 113.700 ;
        RECT 28.640 112.700 28.870 113.340 ;
        RECT 28.620 112.340 28.870 112.700 ;
        RECT 36.930 112.700 37.160 113.340 ;
        RECT 37.420 112.700 37.920 112.900 ;
        RECT 36.930 112.400 37.920 112.700 ;
        RECT 36.930 112.340 37.160 112.400 ;
        RECT 28.620 111.900 28.820 112.340 ;
        RECT 30.525 111.900 35.275 111.980 ;
        RECT 28.020 111.750 35.275 111.900 ;
        RECT 28.020 111.700 30.820 111.750 ;
        RECT 27.450 110.040 27.720 110.300 ;
        RECT 6.220 109.600 6.720 109.900 ;
        RECT 7.080 109.600 7.880 109.680 ;
        RECT 6.220 109.450 7.880 109.600 ;
        RECT 6.220 109.400 7.220 109.450 ;
        RECT 8.120 109.200 8.320 110.040 ;
        RECT 8.720 109.600 9.220 109.900 ;
        RECT 9.510 109.600 10.310 109.680 ;
        RECT 8.720 109.450 10.310 109.600 ;
        RECT 8.720 109.400 9.720 109.450 ;
        RECT 10.520 109.200 10.720 110.040 ;
        RECT 11.120 109.600 11.620 109.900 ;
        RECT 11.940 109.600 12.740 109.680 ;
        RECT 11.120 109.450 12.740 109.600 ;
        RECT 11.120 109.400 12.120 109.450 ;
        RECT 12.920 109.200 13.120 110.040 ;
        RECT 13.520 109.600 14.020 109.900 ;
        RECT 14.370 109.600 15.170 109.680 ;
        RECT 13.520 109.450 15.170 109.600 ;
        RECT 13.520 109.400 14.620 109.450 ;
        RECT 15.420 109.200 15.620 110.040 ;
        RECT 15.920 109.600 16.420 109.900 ;
        RECT 16.800 109.600 17.600 109.680 ;
        RECT 17.820 109.600 18.020 110.040 ;
        RECT 15.920 109.400 18.020 109.600 ;
        RECT 18.420 109.600 18.920 109.900 ;
        RECT 19.230 109.600 20.030 109.680 ;
        RECT 18.420 109.450 20.030 109.600 ;
        RECT 18.420 109.400 19.420 109.450 ;
        RECT 20.220 109.200 20.420 110.040 ;
        RECT 20.820 109.600 21.320 109.900 ;
        RECT 21.660 109.600 22.460 109.680 ;
        RECT 20.820 109.450 22.460 109.600 ;
        RECT 20.820 109.400 21.820 109.450 ;
        RECT 22.620 109.200 22.820 110.040 ;
        RECT 23.320 109.600 23.820 109.900 ;
        RECT 24.090 109.600 24.890 109.680 ;
        RECT 23.320 109.450 24.890 109.600 ;
        RECT 23.320 109.400 24.320 109.450 ;
        RECT 25.120 109.200 25.320 110.040 ;
        RECT 25.720 109.600 26.220 109.900 ;
        RECT 26.520 109.600 27.320 109.680 ;
        RECT 25.720 109.450 27.320 109.600 ;
        RECT 25.720 109.400 26.820 109.450 ;
        RECT 27.520 109.200 27.720 110.040 ;
        RECT 28.020 109.900 28.220 111.700 ;
        RECT 30.880 111.400 34.920 111.430 ;
        RECT 38.120 111.400 38.620 111.700 ;
        RECT 30.880 111.200 38.620 111.400 ;
        RECT 28.640 110.400 28.870 111.040 ;
        RECT 28.620 110.040 28.870 110.400 ;
        RECT 36.930 110.300 37.160 111.040 ;
        RECT 37.420 110.300 37.920 110.500 ;
        RECT 36.930 110.040 37.920 110.300 ;
        RECT 28.620 109.900 28.820 110.040 ;
        RECT 28.020 109.600 28.820 109.900 ;
        RECT 37.020 110.000 37.920 110.040 ;
        RECT 30.525 109.600 35.275 109.680 ;
        RECT 28.020 109.450 35.275 109.600 ;
        RECT 28.020 109.400 30.820 109.450 ;
        RECT 37.020 109.200 37.220 110.000 ;
        RECT 8.120 109.000 37.220 109.200 ;
        RECT 2.300 104.310 36.800 104.400 ;
        RECT 2.300 104.200 39.265 104.310 ;
        RECT 2.300 103.700 3.000 104.200 ;
        RECT 6.220 100.665 6.420 104.200 ;
        RECT 6.720 102.140 6.920 104.200 ;
        RECT 7.220 102.575 7.720 103.300 ;
        RECT 7.220 102.400 7.770 102.575 ;
        RECT 7.230 102.345 7.770 102.400 ;
        RECT 6.720 101.800 6.970 102.140 ;
        RECT 6.170 100.400 6.420 100.665 ;
        RECT 6.170 95.975 6.400 100.400 ;
        RECT 6.740 94.140 6.970 101.800 ;
        RECT 8.030 94.400 8.260 102.140 ;
        RECT 8.620 100.665 8.820 104.200 ;
        RECT 12.120 103.500 12.620 104.000 ;
        RECT 9.720 102.575 10.220 103.300 ;
        RECT 9.660 102.400 10.220 102.575 ;
        RECT 12.120 102.600 12.320 103.500 ;
        RECT 12.120 102.530 12.820 102.600 ;
        RECT 12.120 102.400 13.170 102.530 ;
        RECT 9.660 102.345 10.200 102.400 ;
        RECT 12.120 102.140 12.320 102.400 ;
        RECT 12.630 102.300 13.170 102.400 ;
        RECT 8.600 95.975 8.830 100.665 ;
        RECT 9.170 94.400 9.400 102.140 ;
        RECT 8.030 94.200 9.400 94.400 ;
        RECT 8.030 94.140 8.260 94.200 ;
        RECT 9.170 94.140 9.400 94.200 ;
        RECT 10.460 94.400 10.690 102.140 ;
        RECT 12.120 101.900 12.370 102.140 ;
        RECT 11.570 100.600 11.800 100.630 ;
        RECT 11.570 100.400 11.820 100.600 ;
        RECT 11.570 95.960 11.800 100.400 ;
        RECT 12.140 94.400 12.370 101.900 ;
        RECT 10.460 94.200 12.370 94.400 ;
        RECT 10.460 94.140 10.690 94.200 ;
        RECT 12.140 94.140 12.370 94.200 ;
        RECT 13.430 94.400 13.660 102.140 ;
        RECT 14.520 100.665 14.720 104.200 ;
        RECT 15.120 102.140 15.320 104.200 ;
        RECT 15.620 102.575 16.120 103.300 ;
        RECT 15.620 102.400 16.170 102.575 ;
        RECT 15.630 102.345 16.170 102.400 ;
        RECT 15.120 101.800 15.370 102.140 ;
        RECT 14.520 100.400 14.800 100.665 ;
        RECT 14.570 95.975 14.800 100.400 ;
        RECT 13.430 94.140 13.720 94.400 ;
        RECT 15.140 94.140 15.370 101.800 ;
        RECT 16.430 94.400 16.660 102.140 ;
        RECT 17.020 100.670 17.220 104.200 ;
        RECT 20.820 103.500 21.320 104.000 ;
        RECT 18.020 102.600 18.520 103.300 ;
        RECT 18.020 102.400 20.720 102.600 ;
        RECT 21.020 102.545 21.320 103.500 ;
        RECT 21.020 102.400 21.580 102.545 ;
        RECT 18.060 102.350 18.600 102.400 ;
        RECT 20.520 102.155 20.720 102.400 ;
        RECT 21.040 102.315 21.580 102.400 ;
        RECT 17.000 95.980 17.230 100.670 ;
        RECT 17.570 94.400 17.800 102.145 ;
        RECT 16.430 94.200 17.800 94.400 ;
        RECT 16.430 94.140 16.660 94.200 ;
        RECT 17.570 94.145 17.800 94.200 ;
        RECT 18.860 94.400 19.090 102.145 ;
        RECT 20.520 101.900 20.780 102.155 ;
        RECT 19.980 95.975 20.210 100.645 ;
        RECT 20.550 94.400 20.780 101.900 ;
        RECT 18.860 94.200 20.780 94.400 ;
        RECT 18.860 94.145 19.090 94.200 ;
        RECT 20.550 94.155 20.780 94.200 ;
        RECT 21.840 94.400 22.070 102.155 ;
        RECT 22.920 100.665 23.120 104.200 ;
        RECT 23.520 102.140 23.720 104.200 ;
        RECT 24.020 102.575 24.520 103.300 ;
        RECT 24.020 102.400 24.570 102.575 ;
        RECT 24.030 102.345 24.570 102.400 ;
        RECT 23.520 101.800 23.770 102.140 ;
        RECT 22.920 100.400 23.200 100.665 ;
        RECT 22.970 95.975 23.200 100.400 ;
        RECT 21.840 94.155 22.120 94.400 ;
        RECT 13.520 94.100 13.720 94.140 ;
        RECT 13.520 93.900 14.520 94.100 ;
        RECT 13.620 93.400 14.120 93.700 ;
        RECT 14.320 93.600 14.520 93.900 ;
        RECT 14.320 93.400 16.620 93.600 ;
        RECT 6.620 93.200 14.120 93.400 ;
        RECT 6.620 92.040 6.820 93.200 ;
        RECT 7.220 92.430 7.720 93.000 ;
        RECT 7.210 92.200 7.750 92.430 ;
        RECT 9.120 92.040 9.320 93.200 ;
        RECT 9.620 92.430 10.120 93.000 ;
        RECT 9.620 92.300 10.180 92.430 ;
        RECT 9.640 92.200 10.180 92.300 ;
        RECT 11.520 92.040 11.720 93.200 ;
        RECT 12.020 92.430 12.520 93.000 ;
        RECT 12.020 92.300 12.610 92.430 ;
        RECT 12.070 92.200 12.610 92.300 ;
        RECT 13.920 92.040 14.120 93.200 ;
        RECT 16.420 93.000 16.620 93.400 ;
        RECT 18.520 93.400 19.020 93.700 ;
        RECT 21.920 93.400 22.120 94.155 ;
        RECT 23.540 94.140 23.770 101.800 ;
        RECT 24.830 94.500 25.060 102.140 ;
        RECT 25.320 100.665 25.520 104.200 ;
        RECT 26.420 102.575 26.920 103.300 ;
        RECT 26.420 102.400 26.970 102.575 ;
        RECT 26.430 102.345 26.970 102.400 ;
        RECT 25.320 100.400 25.600 100.665 ;
        RECT 25.370 95.975 25.600 100.400 ;
        RECT 25.940 94.500 26.170 102.140 ;
        RECT 24.830 94.300 26.170 94.500 ;
        RECT 24.830 94.140 25.060 94.300 ;
        RECT 25.940 94.140 26.170 94.300 ;
        RECT 27.230 94.400 27.460 102.140 ;
        RECT 27.720 100.665 27.920 104.200 ;
        RECT 28.320 102.140 28.520 104.200 ;
        RECT 28.820 102.575 29.320 103.300 ;
        RECT 28.820 102.400 29.370 102.575 ;
        RECT 28.830 102.345 29.370 102.400 ;
        RECT 28.320 101.800 28.570 102.140 ;
        RECT 27.720 100.400 28.000 100.665 ;
        RECT 27.770 95.975 28.000 100.400 ;
        RECT 27.230 94.140 27.520 94.400 ;
        RECT 28.340 94.140 28.570 101.800 ;
        RECT 29.630 94.400 29.860 102.140 ;
        RECT 30.120 100.665 30.320 104.200 ;
        RECT 31.920 103.500 32.420 104.000 ;
        RECT 31.220 102.575 31.720 103.300 ;
        RECT 31.220 102.400 31.765 102.575 ;
        RECT 31.225 102.345 31.765 102.400 ;
        RECT 32.120 102.140 32.320 103.500 ;
        RECT 30.120 100.400 30.395 100.665 ;
        RECT 30.165 95.975 30.395 100.400 ;
        RECT 30.735 94.400 30.965 102.140 ;
        RECT 29.630 94.200 30.965 94.400 ;
        RECT 29.630 94.140 29.860 94.200 ;
        RECT 30.735 94.140 30.965 94.200 ;
        RECT 32.025 101.900 32.320 102.140 ;
        RECT 32.025 94.140 32.255 101.900 ;
        RECT 32.620 97.980 32.820 104.200 ;
        RECT 36.575 104.080 39.265 104.200 ;
        RECT 33.400 103.800 33.900 104.000 ;
        RECT 33.400 103.740 36.000 103.800 ;
        RECT 33.400 103.600 39.740 103.740 ;
        RECT 33.400 103.500 33.900 103.600 ;
        RECT 35.740 103.510 39.740 103.600 ;
        RECT 39.945 103.300 40.175 103.460 ;
        RECT 40.900 103.300 41.600 103.800 ;
        RECT 33.420 102.800 33.920 103.300 ;
        RECT 39.945 103.100 41.600 103.300 ;
        RECT 41.900 103.100 42.600 103.800 ;
        RECT 39.945 103.000 40.175 103.100 ;
        RECT 33.170 99.700 33.400 100.245 ;
        RECT 33.120 99.365 33.400 99.700 ;
        RECT 33.720 99.860 33.920 102.800 ;
        RECT 35.740 102.800 39.740 102.950 ;
        RECT 43.900 102.800 44.100 128.600 ;
        RECT 60.975 126.500 65.665 126.550 ;
        RECT 71.000 126.500 73.000 168.300 ;
        RECT 48.400 126.000 48.900 126.500 ;
        RECT 60.975 126.320 73.000 126.500 ;
        RECT 65.400 126.300 73.000 126.320 ;
        RECT 56.800 126.000 58.400 126.100 ;
        RECT 69.200 126.000 69.400 126.300 ;
        RECT 48.400 125.640 48.600 126.000 ;
        RECT 49.040 125.900 58.400 126.000 ;
        RECT 66.800 125.980 69.400 126.000 ;
        RECT 49.040 125.770 57.040 125.900 ;
        RECT 48.400 125.500 48.680 125.640 ;
        RECT 48.450 124.840 48.680 125.500 ;
        RECT 57.200 125.500 57.430 125.510 ;
        RECT 57.200 125.000 58.000 125.500 ;
        RECT 57.200 124.970 57.430 125.000 ;
        RECT 49.040 124.600 57.040 124.710 ;
        RECT 35.740 102.720 44.100 102.800 ;
        RECT 39.400 102.600 44.100 102.720 ;
        RECT 38.020 100.500 38.520 101.000 ;
        RECT 38.020 100.250 38.220 100.500 ;
        RECT 35.980 100.020 40.020 100.250 ;
        RECT 33.720 99.600 33.970 99.860 ;
        RECT 42.030 99.700 42.260 99.860 ;
        RECT 33.740 99.440 33.970 99.600 ;
        RECT 42.020 99.440 42.260 99.700 ;
        RECT 33.120 98.900 33.320 99.365 ;
        RECT 42.020 98.900 42.220 99.440 ;
        RECT 33.120 98.700 43.720 98.900 ;
        RECT 39.220 97.995 43.320 98.000 ;
        RECT 32.620 97.500 32.900 97.980 ;
        RECT 35.480 97.800 43.320 97.995 ;
        RECT 35.480 97.765 39.520 97.800 ;
        RECT 33.240 97.500 33.470 97.560 ;
        RECT 32.620 97.300 33.470 97.500 ;
        RECT 41.530 97.400 41.760 97.560 ;
        RECT 32.670 97.080 32.900 97.300 ;
        RECT 33.240 97.140 33.470 97.300 ;
        RECT 41.520 97.200 42.920 97.400 ;
        RECT 41.530 97.140 41.760 97.200 ;
        RECT 42.720 96.000 42.920 97.200 ;
        RECT 42.420 95.700 42.920 96.000 ;
        RECT 41.420 95.640 42.920 95.700 ;
        RECT 33.760 95.500 42.920 95.640 ;
        RECT 33.760 95.410 41.760 95.500 ;
        RECT 33.170 94.800 33.400 95.280 ;
        RECT 41.920 95.100 42.150 95.150 ;
        RECT 43.120 95.100 43.320 97.800 ;
        RECT 41.920 94.900 43.320 95.100 ;
        RECT 33.170 94.480 33.420 94.800 ;
        RECT 41.920 94.610 42.150 94.900 ;
        RECT 42.420 94.600 42.920 94.900 ;
        RECT 27.320 93.400 27.520 94.140 ;
        RECT 33.220 93.800 33.420 94.480 ;
        RECT 33.760 94.120 41.760 94.350 ;
        RECT 33.820 93.800 34.020 94.120 ;
        RECT 43.520 93.800 43.720 98.700 ;
        RECT 33.220 93.600 43.720 93.800 ;
        RECT 18.520 93.200 26.320 93.400 ;
        RECT 27.320 93.200 42.220 93.400 ;
        RECT 14.520 92.430 15.020 93.000 ;
        RECT 16.420 92.800 17.420 93.000 ;
        RECT 14.500 92.200 15.040 92.430 ;
        RECT 16.420 92.040 16.620 92.800 ;
        RECT 16.920 92.430 17.420 92.800 ;
        RECT 16.920 92.300 17.470 92.430 ;
        RECT 16.930 92.200 17.470 92.300 ;
        RECT 18.820 92.040 19.020 93.200 ;
        RECT 19.420 92.430 19.920 93.000 ;
        RECT 19.360 92.300 19.920 92.430 ;
        RECT 19.360 92.200 19.900 92.300 ;
        RECT 21.220 92.040 21.420 93.200 ;
        RECT 21.820 92.430 22.320 93.000 ;
        RECT 21.790 92.200 22.330 92.430 ;
        RECT 23.720 92.040 23.920 93.200 ;
        RECT 24.220 92.430 24.720 93.000 ;
        RECT 24.220 92.200 24.760 92.430 ;
        RECT 26.120 92.040 26.320 93.200 ;
        RECT 26.620 92.430 27.120 93.000 ;
        RECT 26.620 92.300 27.190 92.430 ;
        RECT 26.650 92.200 27.190 92.300 ;
        RECT 32.155 92.300 38.745 92.330 ;
        RECT 42.020 92.300 42.220 93.200 ;
        RECT 32.155 92.100 42.220 92.300 ;
        RECT 6.620 91.800 6.950 92.040 ;
        RECT 6.720 84.040 6.950 91.800 ;
        RECT 8.010 84.300 8.240 92.040 ;
        RECT 9.120 91.800 9.380 92.040 ;
        RECT 8.010 84.040 8.320 84.300 ;
        RECT 9.150 84.040 9.380 91.800 ;
        RECT 10.440 84.300 10.670 92.040 ;
        RECT 11.520 91.800 11.810 92.040 ;
        RECT 10.440 84.040 10.720 84.300 ;
        RECT 11.580 84.040 11.810 91.800 ;
        RECT 12.870 84.300 13.100 92.040 ;
        RECT 13.920 91.800 14.240 92.040 ;
        RECT 12.870 84.040 13.120 84.300 ;
        RECT 14.010 84.040 14.240 91.800 ;
        RECT 15.300 84.300 15.530 92.040 ;
        RECT 16.420 91.800 16.670 92.040 ;
        RECT 15.300 84.040 15.620 84.300 ;
        RECT 16.440 84.040 16.670 91.800 ;
        RECT 17.730 84.300 17.960 92.040 ;
        RECT 18.820 91.800 19.100 92.040 ;
        RECT 17.730 84.040 18.020 84.300 ;
        RECT 18.870 84.040 19.100 91.800 ;
        RECT 20.160 84.300 20.390 92.040 ;
        RECT 21.220 91.800 21.530 92.040 ;
        RECT 20.160 84.040 20.420 84.300 ;
        RECT 21.300 84.040 21.530 91.800 ;
        RECT 22.590 84.040 22.820 92.040 ;
        RECT 23.720 91.800 23.960 92.040 ;
        RECT 23.730 84.040 23.960 91.800 ;
        RECT 25.020 84.300 25.250 92.040 ;
        RECT 26.120 91.800 26.390 92.040 ;
        RECT 25.020 84.040 25.320 84.300 ;
        RECT 26.160 84.040 26.390 91.800 ;
        RECT 27.450 84.300 27.680 92.040 ;
        RECT 42.020 91.940 42.220 92.100 ;
        RECT 28.640 91.200 28.870 91.940 ;
        RECT 42.020 91.600 42.260 91.940 ;
        RECT 28.620 90.940 28.870 91.200 ;
        RECT 42.030 91.200 42.260 91.600 ;
        RECT 42.520 91.200 43.020 91.500 ;
        RECT 42.030 91.000 43.020 91.200 ;
        RECT 42.030 90.940 42.260 91.000 ;
        RECT 28.620 89.640 28.820 90.940 ;
        RECT 31.800 90.350 39.100 90.580 ;
        RECT 30.880 90.000 34.920 90.030 ;
        RECT 38.120 90.000 38.620 90.200 ;
        RECT 30.880 89.800 38.620 90.000 ;
        RECT 38.120 89.700 38.620 89.800 ;
        RECT 38.820 89.800 39.020 90.350 ;
        RECT 43.220 89.800 43.420 93.600 ;
        RECT 28.620 89.300 28.870 89.640 ;
        RECT 28.640 88.640 28.870 89.300 ;
        RECT 36.930 89.000 37.160 89.640 ;
        RECT 38.820 89.600 43.420 89.800 ;
        RECT 37.420 89.000 37.920 89.200 ;
        RECT 36.930 88.700 37.920 89.000 ;
        RECT 36.930 88.640 37.160 88.700 ;
        RECT 38.820 88.500 39.020 89.600 ;
        RECT 37.420 88.300 39.020 88.500 ;
        RECT 43.900 88.800 44.100 102.600 ;
        RECT 48.000 124.480 57.040 124.600 ;
        RECT 48.000 124.400 49.300 124.480 ;
        RECT 48.000 122.200 48.200 124.400 ;
        RECT 48.400 123.500 48.900 124.000 ;
        RECT 58.200 123.600 58.400 125.900 ;
        RECT 59.140 125.800 69.400 125.980 ;
        RECT 59.140 125.750 67.140 125.800 ;
        RECT 67.400 125.490 68.300 125.500 ;
        RECT 67.345 125.000 68.300 125.490 ;
        RECT 67.345 124.950 67.575 125.000 ;
        RECT 59.140 124.460 67.140 124.690 ;
        RECT 56.800 123.570 58.400 123.600 ;
        RECT 48.400 123.210 48.600 123.500 ;
        RECT 49.040 123.400 58.400 123.570 ;
        RECT 59.200 123.550 59.400 124.460 ;
        RECT 60.975 124.100 65.665 124.120 ;
        RECT 69.200 124.100 69.400 125.800 ;
        RECT 60.975 123.900 69.400 124.100 ;
        RECT 60.975 123.890 65.665 123.900 ;
        RECT 49.040 123.340 57.040 123.400 ;
        RECT 48.400 123.000 48.680 123.210 ;
        RECT 57.300 123.080 58.000 123.100 ;
        RECT 48.450 122.410 48.680 123.000 ;
        RECT 57.200 122.600 58.000 123.080 ;
        RECT 57.200 122.540 57.430 122.600 ;
        RECT 49.040 122.200 57.040 122.280 ;
        RECT 48.000 122.050 57.040 122.200 ;
        RECT 48.000 122.000 49.300 122.050 ;
        RECT 48.000 119.800 48.200 122.000 ;
        RECT 48.400 121.100 48.900 121.600 ;
        RECT 58.200 121.200 58.400 123.400 ;
        RECT 59.140 123.320 67.140 123.550 ;
        RECT 67.345 123.000 67.575 123.060 ;
        RECT 67.345 122.520 68.300 123.000 ;
        RECT 67.400 122.500 68.300 122.520 ;
        RECT 59.140 122.030 67.140 122.260 ;
        RECT 56.800 121.140 58.400 121.200 ;
        RECT 48.400 120.780 48.600 121.100 ;
        RECT 49.040 121.000 58.400 121.140 ;
        RECT 49.040 120.910 57.040 121.000 ;
        RECT 48.400 120.600 48.680 120.780 ;
        RECT 57.300 120.650 58.000 120.700 ;
        RECT 48.450 119.980 48.680 120.600 ;
        RECT 57.200 120.200 58.000 120.650 ;
        RECT 57.200 120.110 57.430 120.200 ;
        RECT 49.040 119.800 57.040 119.850 ;
        RECT 48.000 119.620 57.040 119.800 ;
        RECT 48.000 119.600 49.300 119.620 ;
        RECT 48.000 117.300 48.200 119.600 ;
        RECT 48.400 118.700 48.900 119.200 ;
        RECT 58.200 119.100 58.400 121.000 ;
        RECT 59.200 120.580 59.400 122.030 ;
        RECT 60.960 120.920 65.630 121.150 ;
        RECT 65.400 120.900 65.600 120.920 ;
        RECT 66.900 120.580 69.000 120.600 ;
        RECT 59.140 120.400 69.000 120.580 ;
        RECT 59.140 120.350 67.140 120.400 ;
        RECT 67.400 120.090 67.600 120.400 ;
        RECT 68.500 120.100 69.000 120.400 ;
        RECT 67.300 119.900 67.600 120.090 ;
        RECT 67.300 119.550 67.530 119.900 ;
        RECT 59.140 119.200 67.140 119.290 ;
        RECT 58.200 118.800 58.700 119.100 ;
        RECT 56.800 118.710 58.700 118.800 ;
        RECT 48.400 118.350 48.600 118.700 ;
        RECT 49.040 118.600 58.700 118.710 ;
        RECT 58.900 119.060 67.140 119.200 ;
        RECT 58.900 119.000 59.400 119.060 ;
        RECT 49.040 118.480 57.040 118.600 ;
        RECT 58.900 118.400 59.100 119.000 ;
        RECT 48.400 118.100 48.680 118.350 ;
        RECT 48.450 117.550 48.680 118.100 ;
        RECT 57.200 118.200 57.430 118.220 ;
        RECT 58.400 118.200 59.100 118.400 ;
        RECT 69.200 118.200 69.400 123.900 ;
        RECT 57.200 117.700 58.000 118.200 ;
        RECT 57.200 117.680 57.430 117.700 ;
        RECT 49.040 117.300 57.040 117.420 ;
        RECT 48.000 117.190 57.040 117.300 ;
        RECT 48.000 117.100 49.300 117.190 ;
        RECT 48.000 112.500 48.200 117.100 ;
        RECT 48.400 116.300 48.900 116.800 ;
        RECT 58.400 116.300 58.600 118.200 ;
        RECT 65.400 118.150 69.400 118.200 ;
        RECT 60.975 118.000 69.400 118.150 ;
        RECT 60.975 117.920 65.665 118.000 ;
        RECT 69.200 117.600 69.400 118.000 ;
        RECT 66.800 117.580 69.400 117.600 ;
        RECT 59.140 117.400 69.400 117.580 ;
        RECT 59.140 117.350 67.140 117.400 ;
        RECT 67.400 117.090 68.300 117.100 ;
        RECT 67.345 116.600 68.300 117.090 ;
        RECT 67.345 116.550 67.575 116.600 ;
        RECT 48.400 115.920 48.600 116.300 ;
        RECT 56.800 116.280 58.600 116.300 ;
        RECT 49.040 116.100 58.600 116.280 ;
        RECT 49.040 116.050 57.040 116.100 ;
        RECT 48.400 115.120 48.680 115.920 ;
        RECT 57.800 115.800 58.000 116.100 ;
        RECT 59.140 116.060 67.140 116.290 ;
        RECT 57.300 115.790 58.000 115.800 ;
        RECT 57.200 115.300 58.000 115.790 ;
        RECT 57.200 115.250 57.430 115.300 ;
        RECT 59.200 115.150 59.400 116.060 ;
        RECT 60.980 115.700 65.670 115.720 ;
        RECT 69.200 115.700 69.400 117.400 ;
        RECT 60.980 115.500 69.400 115.700 ;
        RECT 60.980 115.490 65.670 115.500 ;
        RECT 48.400 114.900 48.600 115.120 ;
        RECT 49.040 114.900 57.040 114.990 ;
        RECT 59.145 114.920 67.145 115.150 ;
        RECT 48.400 114.760 57.040 114.900 ;
        RECT 48.400 114.700 49.300 114.760 ;
        RECT 67.400 114.660 68.300 114.700 ;
        RECT 48.400 113.800 48.900 114.300 ;
        RECT 67.350 114.200 68.300 114.660 ;
        RECT 58.200 113.900 58.700 114.200 ;
        RECT 67.350 114.120 67.600 114.200 ;
        RECT 56.800 113.850 58.700 113.900 ;
        RECT 48.400 113.490 48.600 113.800 ;
        RECT 49.040 113.700 58.700 113.850 ;
        RECT 49.040 113.620 57.040 113.700 ;
        RECT 48.400 113.300 48.680 113.490 ;
        RECT 48.450 112.690 48.680 113.300 ;
        RECT 57.200 113.300 57.430 113.360 ;
        RECT 57.200 112.820 58.000 113.300 ;
        RECT 57.300 112.800 58.000 112.820 ;
        RECT 49.040 112.500 57.040 112.560 ;
        RECT 48.000 112.330 57.040 112.500 ;
        RECT 48.000 112.300 49.300 112.330 ;
        RECT 48.000 110.100 48.200 112.300 ;
        RECT 48.400 111.400 48.900 111.900 ;
        RECT 58.200 111.500 58.400 113.700 ;
        RECT 59.145 113.630 67.145 113.860 ;
        RECT 59.200 112.170 59.400 113.630 ;
        RECT 60.975 112.510 65.645 112.740 ;
        RECT 67.400 112.200 67.600 114.120 ;
        RECT 66.900 112.170 67.600 112.200 ;
        RECT 59.155 112.000 67.600 112.170 ;
        RECT 59.155 111.940 67.155 112.000 ;
        RECT 68.500 111.700 69.000 111.900 ;
        RECT 67.400 111.680 69.000 111.700 ;
        RECT 56.800 111.420 58.400 111.500 ;
        RECT 48.400 111.060 48.600 111.400 ;
        RECT 49.040 111.300 58.400 111.420 ;
        RECT 49.040 111.190 57.040 111.300 ;
        RECT 48.400 110.900 48.680 111.060 ;
        RECT 48.450 110.260 48.680 110.900 ;
        RECT 57.200 110.900 57.430 110.930 ;
        RECT 57.200 110.400 58.000 110.900 ;
        RECT 58.200 110.800 58.400 111.300 ;
        RECT 67.315 111.400 69.000 111.680 ;
        RECT 67.315 111.140 67.545 111.400 ;
        RECT 59.155 110.800 67.155 110.880 ;
        RECT 58.200 110.650 67.155 110.800 ;
        RECT 58.200 110.600 59.400 110.650 ;
        RECT 57.200 110.390 57.430 110.400 ;
        RECT 49.040 110.100 57.040 110.130 ;
        RECT 48.000 109.900 57.040 110.100 ;
        RECT 48.000 107.600 48.200 109.900 ;
        RECT 48.400 108.900 48.900 109.400 ;
        RECT 58.200 109.000 58.400 110.600 ;
        RECT 69.200 109.800 69.400 115.500 ;
        RECT 65.400 109.750 69.400 109.800 ;
        RECT 60.975 109.600 69.400 109.750 ;
        RECT 60.975 109.520 65.665 109.600 ;
        RECT 69.200 109.200 69.400 109.600 ;
        RECT 66.800 109.180 69.400 109.200 ;
        RECT 56.800 108.990 58.400 109.000 ;
        RECT 48.400 108.630 48.600 108.900 ;
        RECT 49.040 108.800 58.400 108.990 ;
        RECT 59.140 109.000 69.400 109.180 ;
        RECT 59.140 108.950 67.140 109.000 ;
        RECT 49.040 108.760 57.040 108.800 ;
        RECT 48.400 108.400 48.680 108.630 ;
        RECT 48.450 107.830 48.680 108.400 ;
        RECT 57.200 108.000 58.000 108.500 ;
        RECT 57.200 107.960 57.430 108.000 ;
        RECT 49.040 107.600 57.040 107.700 ;
        RECT 48.000 107.470 57.040 107.600 ;
        RECT 48.000 107.400 49.300 107.470 ;
        RECT 48.000 105.200 48.200 107.400 ;
        RECT 48.400 106.500 48.900 107.000 ;
        RECT 58.200 106.600 58.400 108.800 ;
        RECT 67.400 108.690 68.300 108.700 ;
        RECT 67.345 108.200 68.300 108.690 ;
        RECT 67.345 108.150 67.575 108.200 ;
        RECT 59.140 107.660 67.140 107.890 ;
        RECT 59.300 106.780 59.500 107.660 ;
        RECT 69.200 107.400 69.400 109.000 ;
        RECT 65.400 107.350 69.400 107.400 ;
        RECT 60.975 107.200 69.400 107.350 ;
        RECT 60.975 107.120 65.665 107.200 ;
        RECT 56.800 106.560 58.400 106.600 ;
        RECT 48.400 106.200 48.600 106.500 ;
        RECT 49.040 106.400 58.400 106.560 ;
        RECT 59.140 106.550 67.140 106.780 ;
        RECT 49.040 106.330 57.040 106.400 ;
        RECT 67.400 106.290 68.300 106.300 ;
        RECT 48.400 105.900 48.680 106.200 ;
        RECT 57.300 106.070 58.000 106.100 ;
        RECT 48.450 105.400 48.680 105.900 ;
        RECT 57.200 105.600 58.000 106.070 ;
        RECT 67.345 105.800 68.300 106.290 ;
        RECT 67.345 105.750 67.575 105.800 ;
        RECT 57.200 105.530 57.430 105.600 ;
        RECT 59.140 105.400 67.140 105.490 ;
        RECT 49.040 105.200 57.040 105.270 ;
        RECT 48.000 105.040 57.040 105.200 ;
        RECT 58.200 105.260 67.140 105.400 ;
        RECT 58.200 105.200 59.400 105.260 ;
        RECT 48.000 105.000 49.300 105.040 ;
        RECT 48.000 95.700 48.200 105.000 ;
        RECT 48.400 104.500 53.200 104.700 ;
        RECT 48.400 104.100 48.900 104.500 ;
        RECT 50.700 104.100 50.900 104.500 ;
        RECT 48.400 104.080 49.400 104.100 ;
        RECT 50.700 104.080 51.700 104.100 ;
        RECT 48.400 103.900 50.040 104.080 ;
        RECT 48.400 102.195 48.600 103.900 ;
        RECT 49.040 103.850 50.040 103.900 ;
        RECT 50.700 103.900 52.340 104.080 ;
        RECT 50.700 102.195 50.900 103.900 ;
        RECT 51.340 103.850 52.340 103.900 ;
        RECT 53.000 102.195 53.200 104.500 ;
        RECT 54.300 104.080 56.200 104.100 ;
        RECT 53.640 103.900 56.940 104.080 ;
        RECT 53.640 103.850 54.640 103.900 ;
        RECT 55.940 103.850 56.940 103.900 ;
        RECT 48.400 101.900 48.680 102.195 ;
        RECT 50.700 101.900 50.980 102.195 ;
        RECT 53.000 101.900 53.280 102.195 ;
        RECT 48.450 97.445 48.680 101.900 ;
        RECT 50.200 97.800 50.430 101.840 ;
        RECT 49.040 95.700 50.040 95.790 ;
        RECT 48.000 95.560 50.040 95.700 ;
        RECT 48.000 95.500 49.300 95.560 ;
        RECT 49.000 95.300 49.300 95.500 ;
        RECT 49.000 94.800 49.500 95.300 ;
        RECT 50.200 94.600 50.400 97.800 ;
        RECT 50.750 97.445 50.980 101.900 ;
        RECT 52.500 97.800 52.730 101.840 ;
        RECT 51.340 95.560 52.340 95.790 ;
        RECT 51.400 95.300 51.700 95.560 ;
        RECT 51.400 94.800 51.900 95.300 ;
        RECT 52.500 94.600 52.700 97.800 ;
        RECT 53.050 97.700 53.280 101.900 ;
        RECT 54.800 97.800 55.030 101.840 ;
        RECT 53.050 97.445 53.300 97.700 ;
        RECT 53.100 95.300 53.300 97.445 ;
        RECT 53.640 95.560 54.640 95.790 ;
        RECT 53.700 95.300 54.000 95.560 ;
        RECT 53.100 95.100 53.500 95.300 ;
        RECT 50.200 94.100 50.700 94.600 ;
        RECT 52.500 94.100 53.000 94.600 ;
        RECT 53.300 93.900 53.500 95.100 ;
        RECT 53.700 94.800 54.200 95.300 ;
        RECT 54.800 94.600 55.000 97.800 ;
        RECT 54.700 94.100 55.200 94.600 ;
        RECT 55.350 93.900 55.580 100.920 ;
        RECT 53.300 93.700 55.580 93.900 ;
        RECT 54.600 89.500 54.800 93.700 ;
        RECT 55.350 93.620 55.580 93.700 ;
        RECT 57.100 93.975 57.330 100.565 ;
        RECT 57.100 90.700 57.300 93.975 ;
        RECT 58.200 90.700 58.400 105.200 ;
        RECT 69.200 105.000 69.400 107.200 ;
        RECT 65.400 104.950 69.400 105.000 ;
        RECT 60.975 104.800 69.400 104.950 ;
        RECT 60.975 104.720 65.665 104.800 ;
        RECT 69.200 104.400 69.400 104.800 ;
        RECT 66.800 104.380 69.400 104.400 ;
        RECT 59.140 104.200 69.400 104.380 ;
        RECT 59.140 104.150 67.140 104.200 ;
        RECT 67.400 103.890 68.300 103.900 ;
        RECT 67.345 103.400 68.300 103.890 ;
        RECT 67.345 103.350 67.575 103.400 ;
        RECT 59.140 102.860 67.140 103.090 ;
        RECT 59.200 101.985 59.400 102.860 ;
        RECT 69.200 102.600 69.400 104.200 ;
        RECT 65.400 102.555 69.400 102.600 ;
        RECT 60.975 102.400 69.400 102.555 ;
        RECT 60.975 102.325 65.665 102.400 ;
        RECT 59.140 101.755 67.140 101.985 ;
        RECT 67.400 101.495 68.300 101.500 ;
        RECT 67.345 101.000 68.300 101.495 ;
        RECT 67.345 100.955 67.575 101.000 ;
        RECT 59.140 100.600 67.140 100.695 ;
        RECT 68.500 100.600 69.000 100.800 ;
        RECT 59.140 100.465 69.000 100.600 ;
        RECT 66.900 100.400 69.000 100.465 ;
        RECT 68.500 100.300 69.000 100.400 ;
        RECT 69.200 100.100 69.400 102.400 ;
        RECT 62.300 100.050 69.400 100.100 ;
        RECT 62.080 99.900 69.400 100.050 ;
        RECT 62.080 99.820 62.980 99.900 ;
        RECT 59.480 99.500 60.280 99.550 ;
        RECT 56.600 90.690 58.400 90.700 ;
        RECT 55.940 90.500 58.400 90.690 ;
        RECT 58.600 99.320 60.280 99.500 ;
        RECT 62.300 99.480 62.500 99.820 ;
        RECT 63.700 99.550 64.700 99.600 ;
        RECT 58.600 99.300 59.800 99.320 ;
        RECT 58.600 98.900 58.800 99.300 ;
        RECT 62.140 99.250 62.560 99.480 ;
        RECT 63.700 99.400 65.245 99.550 ;
        RECT 59.120 98.900 59.350 98.960 ;
        RECT 58.600 98.700 59.350 98.900 ;
        RECT 55.940 90.460 56.940 90.500 ;
        RECT 56.000 90.200 56.200 90.460 ;
        RECT 56.000 89.700 56.500 90.200 ;
        RECT 58.600 89.500 58.800 98.700 ;
        RECT 59.120 90.960 59.350 98.700 ;
        RECT 60.410 91.300 60.640 98.960 ;
        RECT 62.765 93.500 62.995 97.240 ;
        RECT 62.765 93.200 63.000 93.500 ;
        RECT 60.410 90.960 60.700 91.300 ;
        RECT 62.200 91.190 62.400 91.200 ;
        RECT 62.140 90.960 62.560 91.190 ;
        RECT 59.610 90.570 60.150 90.800 ;
        RECT 59.900 90.300 60.100 90.570 ;
        RECT 59.600 89.800 60.100 90.300 ;
        RECT 60.500 90.300 60.700 90.960 ;
        RECT 60.500 90.000 61.000 90.300 ;
        RECT 62.200 90.000 62.400 90.960 ;
        RECT 60.500 89.800 62.400 90.000 ;
        RECT 54.600 89.300 58.800 89.500 ;
        RECT 59.900 89.600 60.100 89.800 ;
        RECT 62.800 89.600 63.000 93.200 ;
        RECT 59.900 89.400 63.000 89.600 ;
        RECT 63.700 90.700 63.900 99.400 ;
        RECT 64.365 99.320 65.245 99.400 ;
        RECT 67.800 99.000 68.300 99.300 ;
        RECT 64.600 98.980 68.300 99.000 ;
        RECT 64.440 98.800 68.300 98.980 ;
        RECT 68.500 98.800 69.000 99.300 ;
        RECT 64.440 98.750 64.860 98.800 ;
        RECT 68.600 97.100 68.800 98.800 ;
        RECT 65.020 94.700 65.250 96.740 ;
        RECT 65.020 94.500 66.000 94.700 ;
        RECT 65.020 92.700 65.250 94.500 ;
        RECT 65.500 94.200 66.000 94.500 ;
        RECT 67.720 93.400 67.950 97.100 ;
        RECT 67.600 93.100 67.950 93.400 ;
        RECT 68.510 96.800 68.800 97.100 ;
        RECT 68.510 93.100 68.740 96.800 ;
        RECT 69.200 96.265 69.400 99.900 ;
        RECT 69.080 96.000 69.400 96.265 ;
        RECT 69.080 93.575 69.310 96.000 ;
        RECT 63.700 90.690 64.700 90.700 ;
        RECT 63.700 90.500 64.860 90.690 ;
        RECT 58.600 89.200 58.800 89.300 ;
        RECT 63.700 89.200 63.900 90.500 ;
        RECT 64.440 90.460 64.860 90.500 ;
        RECT 58.600 89.000 63.900 89.200 ;
        RECT 67.600 88.800 67.800 93.100 ;
        RECT 68.000 92.665 68.460 92.895 ;
        RECT 68.100 91.900 68.300 92.665 ;
        RECT 68.100 91.200 68.800 91.900 ;
        RECT 68.100 90.200 68.800 90.900 ;
        RECT 43.900 88.600 67.800 88.800 ;
        RECT 35.020 88.280 37.620 88.300 ;
        RECT 30.525 88.200 37.620 88.280 ;
        RECT 28.020 88.100 37.620 88.200 ;
        RECT 28.020 88.050 35.275 88.100 ;
        RECT 28.020 88.000 30.820 88.050 ;
        RECT 28.020 85.900 28.220 88.000 ;
        RECT 30.880 87.700 34.920 87.730 ;
        RECT 38.120 87.700 38.620 88.000 ;
        RECT 30.880 87.500 38.620 87.700 ;
        RECT 28.640 86.700 28.870 87.340 ;
        RECT 28.620 86.340 28.870 86.700 ;
        RECT 36.930 86.700 37.160 87.340 ;
        RECT 37.420 86.700 37.920 86.900 ;
        RECT 36.930 86.400 37.920 86.700 ;
        RECT 36.930 86.340 37.160 86.400 ;
        RECT 28.620 85.900 28.820 86.340 ;
        RECT 30.525 85.900 35.275 85.980 ;
        RECT 28.020 85.750 35.275 85.900 ;
        RECT 28.020 85.700 30.820 85.750 ;
        RECT 27.450 84.040 27.720 84.300 ;
        RECT 6.220 83.600 6.720 83.900 ;
        RECT 7.080 83.600 7.880 83.680 ;
        RECT 6.220 83.450 7.880 83.600 ;
        RECT 6.220 83.400 7.220 83.450 ;
        RECT 8.120 83.200 8.320 84.040 ;
        RECT 8.720 83.600 9.220 83.900 ;
        RECT 9.510 83.600 10.310 83.680 ;
        RECT 8.720 83.450 10.310 83.600 ;
        RECT 8.720 83.400 9.720 83.450 ;
        RECT 10.520 83.200 10.720 84.040 ;
        RECT 11.120 83.600 11.620 83.900 ;
        RECT 11.940 83.600 12.740 83.680 ;
        RECT 11.120 83.450 12.740 83.600 ;
        RECT 11.120 83.400 12.120 83.450 ;
        RECT 12.920 83.200 13.120 84.040 ;
        RECT 13.520 83.600 14.020 83.900 ;
        RECT 14.370 83.600 15.170 83.680 ;
        RECT 13.520 83.450 15.170 83.600 ;
        RECT 13.520 83.400 14.620 83.450 ;
        RECT 15.420 83.200 15.620 84.040 ;
        RECT 15.920 83.600 16.420 83.900 ;
        RECT 16.800 83.600 17.600 83.680 ;
        RECT 17.820 83.600 18.020 84.040 ;
        RECT 15.920 83.400 18.020 83.600 ;
        RECT 18.420 83.600 18.920 83.900 ;
        RECT 19.230 83.600 20.030 83.680 ;
        RECT 18.420 83.450 20.030 83.600 ;
        RECT 18.420 83.400 19.420 83.450 ;
        RECT 20.220 83.200 20.420 84.040 ;
        RECT 20.820 83.600 21.320 83.900 ;
        RECT 21.660 83.600 22.460 83.680 ;
        RECT 20.820 83.450 22.460 83.600 ;
        RECT 20.820 83.400 21.820 83.450 ;
        RECT 22.620 83.200 22.820 84.040 ;
        RECT 23.320 83.600 23.820 83.900 ;
        RECT 24.090 83.600 24.890 83.680 ;
        RECT 23.320 83.450 24.890 83.600 ;
        RECT 23.320 83.400 24.320 83.450 ;
        RECT 25.120 83.200 25.320 84.040 ;
        RECT 25.720 83.600 26.220 83.900 ;
        RECT 26.520 83.600 27.320 83.680 ;
        RECT 25.720 83.450 27.320 83.600 ;
        RECT 25.720 83.400 26.820 83.450 ;
        RECT 27.520 83.200 27.720 84.040 ;
        RECT 28.020 83.900 28.220 85.700 ;
        RECT 30.880 85.400 34.920 85.430 ;
        RECT 38.120 85.400 38.620 85.700 ;
        RECT 30.880 85.200 38.620 85.400 ;
        RECT 28.640 84.400 28.870 85.040 ;
        RECT 28.620 84.040 28.870 84.400 ;
        RECT 36.930 84.300 37.160 85.040 ;
        RECT 37.420 84.300 37.920 84.500 ;
        RECT 36.930 84.040 37.920 84.300 ;
        RECT 28.620 83.900 28.820 84.040 ;
        RECT 28.020 83.600 28.820 83.900 ;
        RECT 37.020 84.000 37.920 84.040 ;
        RECT 30.525 83.600 35.275 83.680 ;
        RECT 28.020 83.450 35.275 83.600 ;
        RECT 28.020 83.400 30.820 83.450 ;
        RECT 37.020 83.200 37.220 84.000 ;
        RECT 8.120 83.000 37.220 83.200 ;
        RECT 2.300 78.310 36.900 78.400 ;
        RECT 2.300 78.200 39.265 78.310 ;
        RECT 2.300 77.700 3.000 78.200 ;
        RECT 6.220 74.665 6.420 78.200 ;
        RECT 6.720 76.140 6.920 78.200 ;
        RECT 7.220 76.575 7.720 77.300 ;
        RECT 7.220 76.400 7.770 76.575 ;
        RECT 7.230 76.345 7.770 76.400 ;
        RECT 6.720 75.800 6.970 76.140 ;
        RECT 6.170 74.400 6.420 74.665 ;
        RECT 6.170 69.975 6.400 74.400 ;
        RECT 6.740 68.140 6.970 75.800 ;
        RECT 8.030 68.400 8.260 76.140 ;
        RECT 8.620 74.665 8.820 78.200 ;
        RECT 12.120 77.500 12.620 78.000 ;
        RECT 9.720 76.575 10.220 77.300 ;
        RECT 9.660 76.400 10.220 76.575 ;
        RECT 12.120 76.600 12.320 77.500 ;
        RECT 12.120 76.530 12.820 76.600 ;
        RECT 12.120 76.400 13.170 76.530 ;
        RECT 9.660 76.345 10.200 76.400 ;
        RECT 12.120 76.140 12.320 76.400 ;
        RECT 12.630 76.300 13.170 76.400 ;
        RECT 8.600 69.975 8.830 74.665 ;
        RECT 9.170 68.400 9.400 76.140 ;
        RECT 8.030 68.200 9.400 68.400 ;
        RECT 8.030 68.140 8.260 68.200 ;
        RECT 9.170 68.140 9.400 68.200 ;
        RECT 10.460 68.400 10.690 76.140 ;
        RECT 12.120 75.900 12.370 76.140 ;
        RECT 11.570 74.600 11.800 74.630 ;
        RECT 11.570 74.400 11.820 74.600 ;
        RECT 11.570 69.960 11.800 74.400 ;
        RECT 12.140 68.400 12.370 75.900 ;
        RECT 10.460 68.200 12.370 68.400 ;
        RECT 10.460 68.140 10.690 68.200 ;
        RECT 12.140 68.140 12.370 68.200 ;
        RECT 13.430 68.400 13.660 76.140 ;
        RECT 14.520 74.665 14.720 78.200 ;
        RECT 15.120 76.140 15.320 78.200 ;
        RECT 15.620 76.575 16.120 77.300 ;
        RECT 15.620 76.400 16.170 76.575 ;
        RECT 15.630 76.345 16.170 76.400 ;
        RECT 15.120 75.800 15.370 76.140 ;
        RECT 14.520 74.400 14.800 74.665 ;
        RECT 14.570 69.975 14.800 74.400 ;
        RECT 13.430 68.140 13.720 68.400 ;
        RECT 15.140 68.140 15.370 75.800 ;
        RECT 16.430 68.400 16.660 76.140 ;
        RECT 17.020 74.670 17.220 78.200 ;
        RECT 20.820 77.500 21.320 78.000 ;
        RECT 18.020 76.600 18.520 77.300 ;
        RECT 18.020 76.400 20.720 76.600 ;
        RECT 21.020 76.545 21.320 77.500 ;
        RECT 21.020 76.400 21.580 76.545 ;
        RECT 18.060 76.350 18.600 76.400 ;
        RECT 20.520 76.155 20.720 76.400 ;
        RECT 21.040 76.315 21.580 76.400 ;
        RECT 17.000 69.980 17.230 74.670 ;
        RECT 17.570 68.400 17.800 76.145 ;
        RECT 16.430 68.200 17.800 68.400 ;
        RECT 16.430 68.140 16.660 68.200 ;
        RECT 17.570 68.145 17.800 68.200 ;
        RECT 18.860 68.400 19.090 76.145 ;
        RECT 20.520 75.900 20.780 76.155 ;
        RECT 19.980 69.975 20.210 74.645 ;
        RECT 20.550 68.400 20.780 75.900 ;
        RECT 18.860 68.200 20.780 68.400 ;
        RECT 18.860 68.145 19.090 68.200 ;
        RECT 20.550 68.155 20.780 68.200 ;
        RECT 21.840 68.400 22.070 76.155 ;
        RECT 22.920 74.665 23.120 78.200 ;
        RECT 23.520 76.140 23.720 78.200 ;
        RECT 24.020 76.575 24.520 77.300 ;
        RECT 24.020 76.400 24.570 76.575 ;
        RECT 24.030 76.345 24.570 76.400 ;
        RECT 23.520 75.800 23.770 76.140 ;
        RECT 22.920 74.400 23.200 74.665 ;
        RECT 22.970 69.975 23.200 74.400 ;
        RECT 21.840 68.155 22.120 68.400 ;
        RECT 13.520 68.100 13.720 68.140 ;
        RECT 13.520 67.900 14.520 68.100 ;
        RECT 13.620 67.400 14.120 67.700 ;
        RECT 14.320 67.600 14.520 67.900 ;
        RECT 14.320 67.400 16.620 67.600 ;
        RECT 6.620 67.200 14.120 67.400 ;
        RECT 6.620 66.040 6.820 67.200 ;
        RECT 7.220 66.430 7.720 67.000 ;
        RECT 7.210 66.200 7.750 66.430 ;
        RECT 9.120 66.040 9.320 67.200 ;
        RECT 9.620 66.430 10.120 67.000 ;
        RECT 9.620 66.300 10.180 66.430 ;
        RECT 9.640 66.200 10.180 66.300 ;
        RECT 11.520 66.040 11.720 67.200 ;
        RECT 12.020 66.430 12.520 67.000 ;
        RECT 12.020 66.300 12.610 66.430 ;
        RECT 12.070 66.200 12.610 66.300 ;
        RECT 13.920 66.040 14.120 67.200 ;
        RECT 16.420 67.000 16.620 67.400 ;
        RECT 18.520 67.400 19.020 67.700 ;
        RECT 21.920 67.400 22.120 68.155 ;
        RECT 23.540 68.140 23.770 75.800 ;
        RECT 24.830 68.500 25.060 76.140 ;
        RECT 25.320 74.665 25.520 78.200 ;
        RECT 26.420 76.575 26.920 77.300 ;
        RECT 26.420 76.400 26.970 76.575 ;
        RECT 26.430 76.345 26.970 76.400 ;
        RECT 25.320 74.400 25.600 74.665 ;
        RECT 25.370 69.975 25.600 74.400 ;
        RECT 25.940 68.500 26.170 76.140 ;
        RECT 24.830 68.300 26.170 68.500 ;
        RECT 24.830 68.140 25.060 68.300 ;
        RECT 25.940 68.140 26.170 68.300 ;
        RECT 27.230 68.400 27.460 76.140 ;
        RECT 27.720 74.665 27.920 78.200 ;
        RECT 28.320 76.140 28.520 78.200 ;
        RECT 28.820 76.575 29.320 77.300 ;
        RECT 28.820 76.400 29.370 76.575 ;
        RECT 28.830 76.345 29.370 76.400 ;
        RECT 28.320 75.800 28.570 76.140 ;
        RECT 27.720 74.400 28.000 74.665 ;
        RECT 27.770 69.975 28.000 74.400 ;
        RECT 27.230 68.140 27.520 68.400 ;
        RECT 28.340 68.140 28.570 75.800 ;
        RECT 29.630 68.400 29.860 76.140 ;
        RECT 30.120 74.665 30.320 78.200 ;
        RECT 31.920 77.500 32.420 78.000 ;
        RECT 31.220 76.575 31.720 77.300 ;
        RECT 31.220 76.400 31.765 76.575 ;
        RECT 31.225 76.345 31.765 76.400 ;
        RECT 32.120 76.140 32.320 77.500 ;
        RECT 30.120 74.400 30.395 74.665 ;
        RECT 30.165 69.975 30.395 74.400 ;
        RECT 30.735 68.400 30.965 76.140 ;
        RECT 29.630 68.200 30.965 68.400 ;
        RECT 29.630 68.140 29.860 68.200 ;
        RECT 30.735 68.140 30.965 68.200 ;
        RECT 32.025 75.900 32.320 76.140 ;
        RECT 32.025 68.140 32.255 75.900 ;
        RECT 32.620 71.980 32.820 78.200 ;
        RECT 36.575 78.080 39.265 78.200 ;
        RECT 33.400 77.800 33.900 78.000 ;
        RECT 33.400 77.740 36.000 77.800 ;
        RECT 33.400 77.600 39.740 77.740 ;
        RECT 33.400 77.500 33.900 77.600 ;
        RECT 35.740 77.510 39.740 77.600 ;
        RECT 39.945 77.300 40.175 77.460 ;
        RECT 40.900 77.300 41.600 77.800 ;
        RECT 33.420 76.800 33.920 77.300 ;
        RECT 39.945 77.100 41.600 77.300 ;
        RECT 41.900 77.100 42.600 77.800 ;
        RECT 39.945 77.000 40.175 77.100 ;
        RECT 33.170 73.700 33.400 74.245 ;
        RECT 33.120 73.365 33.400 73.700 ;
        RECT 33.720 73.860 33.920 76.800 ;
        RECT 35.740 76.800 39.740 76.950 ;
        RECT 43.900 76.800 44.100 88.600 ;
        RECT 60.975 84.500 65.665 84.550 ;
        RECT 71.000 84.500 73.000 126.300 ;
        RECT 48.400 84.000 48.900 84.500 ;
        RECT 60.975 84.320 73.000 84.500 ;
        RECT 65.400 84.300 73.000 84.320 ;
        RECT 56.800 84.000 58.400 84.100 ;
        RECT 69.200 84.000 69.400 84.300 ;
        RECT 48.400 83.640 48.600 84.000 ;
        RECT 49.040 83.900 58.400 84.000 ;
        RECT 66.800 83.980 69.400 84.000 ;
        RECT 49.040 83.770 57.040 83.900 ;
        RECT 48.400 83.500 48.680 83.640 ;
        RECT 48.450 82.840 48.680 83.500 ;
        RECT 57.200 83.500 57.430 83.510 ;
        RECT 57.200 83.000 58.000 83.500 ;
        RECT 57.200 82.970 57.430 83.000 ;
        RECT 49.040 82.600 57.040 82.710 ;
        RECT 35.740 76.720 44.100 76.800 ;
        RECT 39.400 76.600 44.100 76.720 ;
        RECT 38.020 74.500 38.520 75.000 ;
        RECT 38.020 74.250 38.220 74.500 ;
        RECT 35.980 74.020 40.020 74.250 ;
        RECT 33.720 73.600 33.970 73.860 ;
        RECT 42.030 73.700 42.260 73.860 ;
        RECT 33.740 73.440 33.970 73.600 ;
        RECT 42.020 73.440 42.260 73.700 ;
        RECT 33.120 72.900 33.320 73.365 ;
        RECT 42.020 72.900 42.220 73.440 ;
        RECT 33.120 72.700 43.720 72.900 ;
        RECT 39.220 71.995 43.320 72.000 ;
        RECT 32.620 71.500 32.900 71.980 ;
        RECT 35.480 71.800 43.320 71.995 ;
        RECT 35.480 71.765 39.520 71.800 ;
        RECT 33.240 71.500 33.470 71.560 ;
        RECT 32.620 71.300 33.470 71.500 ;
        RECT 41.530 71.400 41.760 71.560 ;
        RECT 32.670 71.080 32.900 71.300 ;
        RECT 33.240 71.140 33.470 71.300 ;
        RECT 41.520 71.200 42.920 71.400 ;
        RECT 41.530 71.140 41.760 71.200 ;
        RECT 42.720 70.000 42.920 71.200 ;
        RECT 42.420 69.700 42.920 70.000 ;
        RECT 41.420 69.640 42.920 69.700 ;
        RECT 33.760 69.500 42.920 69.640 ;
        RECT 33.760 69.410 41.760 69.500 ;
        RECT 33.170 68.800 33.400 69.280 ;
        RECT 41.920 69.100 42.150 69.150 ;
        RECT 43.120 69.100 43.320 71.800 ;
        RECT 41.920 68.900 43.320 69.100 ;
        RECT 33.170 68.480 33.420 68.800 ;
        RECT 41.920 68.610 42.150 68.900 ;
        RECT 42.420 68.600 42.920 68.900 ;
        RECT 27.320 67.400 27.520 68.140 ;
        RECT 33.220 67.800 33.420 68.480 ;
        RECT 33.760 68.120 41.760 68.350 ;
        RECT 33.820 67.800 34.020 68.120 ;
        RECT 43.520 67.800 43.720 72.700 ;
        RECT 33.220 67.600 43.720 67.800 ;
        RECT 18.520 67.200 26.320 67.400 ;
        RECT 27.320 67.200 42.220 67.400 ;
        RECT 14.520 66.430 15.020 67.000 ;
        RECT 16.420 66.800 17.420 67.000 ;
        RECT 14.500 66.200 15.040 66.430 ;
        RECT 16.420 66.040 16.620 66.800 ;
        RECT 16.920 66.430 17.420 66.800 ;
        RECT 16.920 66.300 17.470 66.430 ;
        RECT 16.930 66.200 17.470 66.300 ;
        RECT 18.820 66.040 19.020 67.200 ;
        RECT 19.420 66.430 19.920 67.000 ;
        RECT 19.360 66.300 19.920 66.430 ;
        RECT 19.360 66.200 19.900 66.300 ;
        RECT 21.220 66.040 21.420 67.200 ;
        RECT 21.820 66.430 22.320 67.000 ;
        RECT 21.790 66.200 22.330 66.430 ;
        RECT 23.720 66.040 23.920 67.200 ;
        RECT 24.220 66.430 24.720 67.000 ;
        RECT 24.220 66.200 24.760 66.430 ;
        RECT 26.120 66.040 26.320 67.200 ;
        RECT 26.620 66.430 27.120 67.000 ;
        RECT 26.620 66.300 27.190 66.430 ;
        RECT 26.650 66.200 27.190 66.300 ;
        RECT 32.155 66.300 38.745 66.330 ;
        RECT 42.020 66.300 42.220 67.200 ;
        RECT 32.155 66.100 42.220 66.300 ;
        RECT 6.620 65.800 6.950 66.040 ;
        RECT 6.720 58.040 6.950 65.800 ;
        RECT 8.010 58.300 8.240 66.040 ;
        RECT 9.120 65.800 9.380 66.040 ;
        RECT 8.010 58.040 8.320 58.300 ;
        RECT 9.150 58.040 9.380 65.800 ;
        RECT 10.440 58.300 10.670 66.040 ;
        RECT 11.520 65.800 11.810 66.040 ;
        RECT 10.440 58.040 10.720 58.300 ;
        RECT 11.580 58.040 11.810 65.800 ;
        RECT 12.870 58.300 13.100 66.040 ;
        RECT 13.920 65.800 14.240 66.040 ;
        RECT 12.870 58.040 13.120 58.300 ;
        RECT 14.010 58.040 14.240 65.800 ;
        RECT 15.300 58.300 15.530 66.040 ;
        RECT 16.420 65.800 16.670 66.040 ;
        RECT 15.300 58.040 15.620 58.300 ;
        RECT 16.440 58.040 16.670 65.800 ;
        RECT 17.730 58.300 17.960 66.040 ;
        RECT 18.820 65.800 19.100 66.040 ;
        RECT 17.730 58.040 18.020 58.300 ;
        RECT 18.870 58.040 19.100 65.800 ;
        RECT 20.160 58.300 20.390 66.040 ;
        RECT 21.220 65.800 21.530 66.040 ;
        RECT 20.160 58.040 20.420 58.300 ;
        RECT 21.300 58.040 21.530 65.800 ;
        RECT 22.590 58.040 22.820 66.040 ;
        RECT 23.720 65.800 23.960 66.040 ;
        RECT 23.730 58.040 23.960 65.800 ;
        RECT 25.020 58.300 25.250 66.040 ;
        RECT 26.120 65.800 26.390 66.040 ;
        RECT 25.020 58.040 25.320 58.300 ;
        RECT 26.160 58.040 26.390 65.800 ;
        RECT 27.450 58.300 27.680 66.040 ;
        RECT 42.020 65.940 42.220 66.100 ;
        RECT 28.640 65.200 28.870 65.940 ;
        RECT 42.020 65.600 42.260 65.940 ;
        RECT 28.620 64.940 28.870 65.200 ;
        RECT 42.030 65.200 42.260 65.600 ;
        RECT 42.520 65.200 43.020 65.500 ;
        RECT 42.030 65.000 43.020 65.200 ;
        RECT 42.030 64.940 42.260 65.000 ;
        RECT 28.620 63.640 28.820 64.940 ;
        RECT 31.800 64.350 39.100 64.580 ;
        RECT 30.880 64.000 34.920 64.030 ;
        RECT 38.120 64.000 38.620 64.200 ;
        RECT 30.880 63.800 38.620 64.000 ;
        RECT 38.120 63.700 38.620 63.800 ;
        RECT 38.820 63.800 39.020 64.350 ;
        RECT 43.220 63.800 43.420 67.600 ;
        RECT 28.620 63.300 28.870 63.640 ;
        RECT 28.640 62.640 28.870 63.300 ;
        RECT 36.930 63.000 37.160 63.640 ;
        RECT 38.820 63.600 43.420 63.800 ;
        RECT 37.420 63.000 37.920 63.200 ;
        RECT 36.930 62.700 37.920 63.000 ;
        RECT 36.930 62.640 37.160 62.700 ;
        RECT 38.820 62.500 39.020 63.600 ;
        RECT 37.420 62.300 39.020 62.500 ;
        RECT 35.020 62.280 37.620 62.300 ;
        RECT 30.525 62.200 37.620 62.280 ;
        RECT 28.020 62.100 37.620 62.200 ;
        RECT 28.020 62.050 35.275 62.100 ;
        RECT 28.020 62.000 30.820 62.050 ;
        RECT 28.020 59.900 28.220 62.000 ;
        RECT 30.880 61.700 34.920 61.730 ;
        RECT 38.120 61.700 38.620 62.000 ;
        RECT 30.880 61.500 38.620 61.700 ;
        RECT 28.640 60.700 28.870 61.340 ;
        RECT 28.620 60.340 28.870 60.700 ;
        RECT 36.930 60.700 37.160 61.340 ;
        RECT 37.420 60.700 37.920 60.900 ;
        RECT 36.930 60.400 37.920 60.700 ;
        RECT 36.930 60.340 37.160 60.400 ;
        RECT 28.620 59.900 28.820 60.340 ;
        RECT 30.525 59.900 35.275 59.980 ;
        RECT 28.020 59.750 35.275 59.900 ;
        RECT 28.020 59.700 30.820 59.750 ;
        RECT 27.450 58.040 27.720 58.300 ;
        RECT 6.220 57.600 6.720 57.900 ;
        RECT 7.080 57.600 7.880 57.680 ;
        RECT 6.220 57.450 7.880 57.600 ;
        RECT 6.220 57.400 7.220 57.450 ;
        RECT 8.120 57.200 8.320 58.040 ;
        RECT 8.720 57.600 9.220 57.900 ;
        RECT 9.510 57.600 10.310 57.680 ;
        RECT 8.720 57.450 10.310 57.600 ;
        RECT 8.720 57.400 9.720 57.450 ;
        RECT 10.520 57.200 10.720 58.040 ;
        RECT 11.120 57.600 11.620 57.900 ;
        RECT 11.940 57.600 12.740 57.680 ;
        RECT 11.120 57.450 12.740 57.600 ;
        RECT 11.120 57.400 12.120 57.450 ;
        RECT 12.920 57.200 13.120 58.040 ;
        RECT 13.520 57.600 14.020 57.900 ;
        RECT 14.370 57.600 15.170 57.680 ;
        RECT 13.520 57.450 15.170 57.600 ;
        RECT 13.520 57.400 14.620 57.450 ;
        RECT 15.420 57.200 15.620 58.040 ;
        RECT 15.920 57.600 16.420 57.900 ;
        RECT 16.800 57.600 17.600 57.680 ;
        RECT 17.820 57.600 18.020 58.040 ;
        RECT 15.920 57.400 18.020 57.600 ;
        RECT 18.420 57.600 18.920 57.900 ;
        RECT 19.230 57.600 20.030 57.680 ;
        RECT 18.420 57.450 20.030 57.600 ;
        RECT 18.420 57.400 19.420 57.450 ;
        RECT 20.220 57.200 20.420 58.040 ;
        RECT 20.820 57.600 21.320 57.900 ;
        RECT 21.660 57.600 22.460 57.680 ;
        RECT 20.820 57.450 22.460 57.600 ;
        RECT 20.820 57.400 21.820 57.450 ;
        RECT 22.620 57.200 22.820 58.040 ;
        RECT 23.320 57.600 23.820 57.900 ;
        RECT 24.090 57.600 24.890 57.680 ;
        RECT 23.320 57.450 24.890 57.600 ;
        RECT 23.320 57.400 24.320 57.450 ;
        RECT 25.120 57.200 25.320 58.040 ;
        RECT 25.720 57.600 26.220 57.900 ;
        RECT 26.520 57.600 27.320 57.680 ;
        RECT 25.720 57.450 27.320 57.600 ;
        RECT 25.720 57.400 26.820 57.450 ;
        RECT 27.520 57.200 27.720 58.040 ;
        RECT 28.020 57.900 28.220 59.700 ;
        RECT 30.880 59.400 34.920 59.430 ;
        RECT 38.120 59.400 38.620 59.700 ;
        RECT 30.880 59.200 38.620 59.400 ;
        RECT 28.640 58.400 28.870 59.040 ;
        RECT 28.620 58.040 28.870 58.400 ;
        RECT 36.930 58.300 37.160 59.040 ;
        RECT 37.420 58.300 37.920 58.500 ;
        RECT 36.930 58.040 37.920 58.300 ;
        RECT 28.620 57.900 28.820 58.040 ;
        RECT 28.020 57.600 28.820 57.900 ;
        RECT 37.020 58.000 37.920 58.040 ;
        RECT 30.525 57.600 35.275 57.680 ;
        RECT 28.020 57.450 35.275 57.600 ;
        RECT 28.020 57.400 30.820 57.450 ;
        RECT 37.020 57.200 37.220 58.000 ;
        RECT 8.120 57.000 37.220 57.200 ;
        RECT 2.300 52.310 36.900 52.400 ;
        RECT 2.300 52.200 39.265 52.310 ;
        RECT 2.300 51.700 3.000 52.200 ;
        RECT 6.220 48.665 6.420 52.200 ;
        RECT 6.720 50.140 6.920 52.200 ;
        RECT 7.220 50.575 7.720 51.300 ;
        RECT 7.220 50.400 7.770 50.575 ;
        RECT 7.230 50.345 7.770 50.400 ;
        RECT 6.720 49.800 6.970 50.140 ;
        RECT 6.170 48.400 6.420 48.665 ;
        RECT 6.170 43.975 6.400 48.400 ;
        RECT 6.740 42.140 6.970 49.800 ;
        RECT 8.030 42.400 8.260 50.140 ;
        RECT 8.620 48.665 8.820 52.200 ;
        RECT 12.120 51.500 12.620 52.000 ;
        RECT 9.720 50.575 10.220 51.300 ;
        RECT 9.660 50.400 10.220 50.575 ;
        RECT 12.120 50.600 12.320 51.500 ;
        RECT 12.120 50.530 12.820 50.600 ;
        RECT 12.120 50.400 13.170 50.530 ;
        RECT 9.660 50.345 10.200 50.400 ;
        RECT 12.120 50.140 12.320 50.400 ;
        RECT 12.630 50.300 13.170 50.400 ;
        RECT 8.600 43.975 8.830 48.665 ;
        RECT 9.170 42.400 9.400 50.140 ;
        RECT 8.030 42.200 9.400 42.400 ;
        RECT 8.030 42.140 8.260 42.200 ;
        RECT 9.170 42.140 9.400 42.200 ;
        RECT 10.460 42.400 10.690 50.140 ;
        RECT 12.120 49.900 12.370 50.140 ;
        RECT 11.570 48.600 11.800 48.630 ;
        RECT 11.570 48.400 11.820 48.600 ;
        RECT 11.570 43.960 11.800 48.400 ;
        RECT 12.140 42.400 12.370 49.900 ;
        RECT 10.460 42.200 12.370 42.400 ;
        RECT 10.460 42.140 10.690 42.200 ;
        RECT 12.140 42.140 12.370 42.200 ;
        RECT 13.430 42.400 13.660 50.140 ;
        RECT 14.520 48.665 14.720 52.200 ;
        RECT 15.120 50.140 15.320 52.200 ;
        RECT 15.620 50.575 16.120 51.300 ;
        RECT 15.620 50.400 16.170 50.575 ;
        RECT 15.630 50.345 16.170 50.400 ;
        RECT 15.120 49.800 15.370 50.140 ;
        RECT 14.520 48.400 14.800 48.665 ;
        RECT 14.570 43.975 14.800 48.400 ;
        RECT 13.430 42.140 13.720 42.400 ;
        RECT 15.140 42.140 15.370 49.800 ;
        RECT 16.430 42.400 16.660 50.140 ;
        RECT 17.020 48.670 17.220 52.200 ;
        RECT 20.820 51.500 21.320 52.000 ;
        RECT 18.020 50.600 18.520 51.300 ;
        RECT 18.020 50.400 20.720 50.600 ;
        RECT 21.020 50.545 21.320 51.500 ;
        RECT 21.020 50.400 21.580 50.545 ;
        RECT 18.060 50.350 18.600 50.400 ;
        RECT 20.520 50.155 20.720 50.400 ;
        RECT 21.040 50.315 21.580 50.400 ;
        RECT 17.000 43.980 17.230 48.670 ;
        RECT 17.570 42.400 17.800 50.145 ;
        RECT 16.430 42.200 17.800 42.400 ;
        RECT 16.430 42.140 16.660 42.200 ;
        RECT 17.570 42.145 17.800 42.200 ;
        RECT 18.860 42.400 19.090 50.145 ;
        RECT 20.520 49.900 20.780 50.155 ;
        RECT 19.980 43.975 20.210 48.645 ;
        RECT 20.550 42.400 20.780 49.900 ;
        RECT 18.860 42.200 20.780 42.400 ;
        RECT 18.860 42.145 19.090 42.200 ;
        RECT 20.550 42.155 20.780 42.200 ;
        RECT 21.840 42.400 22.070 50.155 ;
        RECT 22.920 48.665 23.120 52.200 ;
        RECT 23.520 50.140 23.720 52.200 ;
        RECT 24.020 50.575 24.520 51.300 ;
        RECT 24.020 50.400 24.570 50.575 ;
        RECT 24.030 50.345 24.570 50.400 ;
        RECT 23.520 49.800 23.770 50.140 ;
        RECT 22.920 48.400 23.200 48.665 ;
        RECT 22.970 43.975 23.200 48.400 ;
        RECT 21.840 42.155 22.120 42.400 ;
        RECT 13.520 42.100 13.720 42.140 ;
        RECT 13.520 41.900 14.520 42.100 ;
        RECT 13.620 41.400 14.120 41.700 ;
        RECT 14.320 41.600 14.520 41.900 ;
        RECT 14.320 41.400 16.620 41.600 ;
        RECT 6.620 41.200 14.120 41.400 ;
        RECT 6.620 40.040 6.820 41.200 ;
        RECT 7.220 40.430 7.720 41.000 ;
        RECT 7.210 40.200 7.750 40.430 ;
        RECT 9.120 40.040 9.320 41.200 ;
        RECT 9.620 40.430 10.120 41.000 ;
        RECT 9.620 40.300 10.180 40.430 ;
        RECT 9.640 40.200 10.180 40.300 ;
        RECT 11.520 40.040 11.720 41.200 ;
        RECT 12.020 40.430 12.520 41.000 ;
        RECT 12.020 40.300 12.610 40.430 ;
        RECT 12.070 40.200 12.610 40.300 ;
        RECT 13.920 40.040 14.120 41.200 ;
        RECT 16.420 41.000 16.620 41.400 ;
        RECT 18.520 41.400 19.020 41.700 ;
        RECT 21.920 41.400 22.120 42.155 ;
        RECT 23.540 42.140 23.770 49.800 ;
        RECT 24.830 42.500 25.060 50.140 ;
        RECT 25.320 48.665 25.520 52.200 ;
        RECT 26.420 50.575 26.920 51.300 ;
        RECT 26.420 50.400 26.970 50.575 ;
        RECT 26.430 50.345 26.970 50.400 ;
        RECT 25.320 48.400 25.600 48.665 ;
        RECT 25.370 43.975 25.600 48.400 ;
        RECT 25.940 42.500 26.170 50.140 ;
        RECT 24.830 42.300 26.170 42.500 ;
        RECT 24.830 42.140 25.060 42.300 ;
        RECT 25.940 42.140 26.170 42.300 ;
        RECT 27.230 42.400 27.460 50.140 ;
        RECT 27.720 48.665 27.920 52.200 ;
        RECT 28.320 50.140 28.520 52.200 ;
        RECT 28.820 50.575 29.320 51.300 ;
        RECT 28.820 50.400 29.370 50.575 ;
        RECT 28.830 50.345 29.370 50.400 ;
        RECT 28.320 49.800 28.570 50.140 ;
        RECT 27.720 48.400 28.000 48.665 ;
        RECT 27.770 43.975 28.000 48.400 ;
        RECT 27.230 42.140 27.520 42.400 ;
        RECT 28.340 42.140 28.570 49.800 ;
        RECT 29.630 42.400 29.860 50.140 ;
        RECT 30.120 48.665 30.320 52.200 ;
        RECT 31.920 51.500 32.420 52.000 ;
        RECT 31.220 50.575 31.720 51.300 ;
        RECT 31.220 50.400 31.765 50.575 ;
        RECT 31.225 50.345 31.765 50.400 ;
        RECT 32.120 50.140 32.320 51.500 ;
        RECT 30.120 48.400 30.395 48.665 ;
        RECT 30.165 43.975 30.395 48.400 ;
        RECT 30.735 42.400 30.965 50.140 ;
        RECT 29.630 42.200 30.965 42.400 ;
        RECT 29.630 42.140 29.860 42.200 ;
        RECT 30.735 42.140 30.965 42.200 ;
        RECT 32.025 49.900 32.320 50.140 ;
        RECT 32.025 42.140 32.255 49.900 ;
        RECT 32.620 45.980 32.820 52.200 ;
        RECT 36.575 52.080 39.265 52.200 ;
        RECT 33.400 51.800 33.900 52.000 ;
        RECT 33.400 51.740 36.100 51.800 ;
        RECT 33.400 51.600 39.740 51.740 ;
        RECT 33.400 51.500 33.900 51.600 ;
        RECT 35.740 51.510 39.740 51.600 ;
        RECT 39.945 51.300 40.175 51.460 ;
        RECT 40.900 51.300 41.600 51.800 ;
        RECT 33.420 50.800 33.920 51.300 ;
        RECT 39.945 51.100 41.600 51.300 ;
        RECT 41.900 51.100 42.600 51.800 ;
        RECT 39.945 51.000 40.175 51.100 ;
        RECT 33.170 47.700 33.400 48.245 ;
        RECT 33.120 47.365 33.400 47.700 ;
        RECT 33.720 47.860 33.920 50.800 ;
        RECT 35.740 50.900 39.740 50.950 ;
        RECT 35.740 50.800 39.800 50.900 ;
        RECT 43.900 50.800 44.100 76.600 ;
        RECT 48.000 82.480 57.040 82.600 ;
        RECT 48.000 82.400 49.300 82.480 ;
        RECT 48.000 80.200 48.200 82.400 ;
        RECT 48.400 81.500 48.900 82.000 ;
        RECT 58.200 81.600 58.400 83.900 ;
        RECT 59.140 83.800 69.400 83.980 ;
        RECT 59.140 83.750 67.140 83.800 ;
        RECT 67.400 83.490 68.300 83.500 ;
        RECT 67.345 83.000 68.300 83.490 ;
        RECT 67.345 82.950 67.575 83.000 ;
        RECT 59.140 82.460 67.140 82.690 ;
        RECT 56.800 81.570 58.400 81.600 ;
        RECT 48.400 81.210 48.600 81.500 ;
        RECT 49.040 81.400 58.400 81.570 ;
        RECT 59.200 81.550 59.400 82.460 ;
        RECT 60.975 82.100 65.665 82.120 ;
        RECT 69.200 82.100 69.400 83.800 ;
        RECT 60.975 81.900 69.400 82.100 ;
        RECT 60.975 81.890 65.665 81.900 ;
        RECT 49.040 81.340 57.040 81.400 ;
        RECT 48.400 81.000 48.680 81.210 ;
        RECT 57.300 81.080 58.000 81.100 ;
        RECT 48.450 80.410 48.680 81.000 ;
        RECT 57.200 80.600 58.000 81.080 ;
        RECT 57.200 80.540 57.430 80.600 ;
        RECT 49.040 80.200 57.040 80.280 ;
        RECT 48.000 80.050 57.040 80.200 ;
        RECT 48.000 80.000 49.300 80.050 ;
        RECT 48.000 77.800 48.200 80.000 ;
        RECT 48.400 79.100 48.900 79.600 ;
        RECT 58.200 79.200 58.400 81.400 ;
        RECT 59.140 81.320 67.140 81.550 ;
        RECT 67.345 81.000 67.575 81.060 ;
        RECT 67.345 80.520 68.300 81.000 ;
        RECT 67.400 80.500 68.300 80.520 ;
        RECT 59.140 80.030 67.140 80.260 ;
        RECT 56.800 79.140 58.400 79.200 ;
        RECT 48.400 78.780 48.600 79.100 ;
        RECT 49.040 79.000 58.400 79.140 ;
        RECT 49.040 78.910 57.040 79.000 ;
        RECT 48.400 78.600 48.680 78.780 ;
        RECT 57.300 78.650 58.000 78.700 ;
        RECT 48.450 77.980 48.680 78.600 ;
        RECT 57.200 78.200 58.000 78.650 ;
        RECT 57.200 78.110 57.430 78.200 ;
        RECT 49.040 77.800 57.040 77.850 ;
        RECT 48.000 77.620 57.040 77.800 ;
        RECT 48.000 77.600 49.300 77.620 ;
        RECT 48.000 75.300 48.200 77.600 ;
        RECT 48.400 76.700 48.900 77.200 ;
        RECT 58.200 77.100 58.400 79.000 ;
        RECT 59.200 78.580 59.400 80.030 ;
        RECT 60.960 78.920 65.630 79.150 ;
        RECT 65.400 78.900 65.600 78.920 ;
        RECT 66.900 78.580 69.000 78.600 ;
        RECT 59.140 78.400 69.000 78.580 ;
        RECT 59.140 78.350 67.140 78.400 ;
        RECT 67.400 78.090 67.600 78.400 ;
        RECT 68.500 78.100 69.000 78.400 ;
        RECT 67.300 77.900 67.600 78.090 ;
        RECT 67.300 77.550 67.530 77.900 ;
        RECT 59.140 77.200 67.140 77.290 ;
        RECT 58.200 76.800 58.700 77.100 ;
        RECT 56.800 76.710 58.700 76.800 ;
        RECT 48.400 76.350 48.600 76.700 ;
        RECT 49.040 76.600 58.700 76.710 ;
        RECT 58.900 77.060 67.140 77.200 ;
        RECT 58.900 77.000 59.400 77.060 ;
        RECT 49.040 76.480 57.040 76.600 ;
        RECT 58.900 76.400 59.100 77.000 ;
        RECT 48.400 76.100 48.680 76.350 ;
        RECT 48.450 75.550 48.680 76.100 ;
        RECT 57.200 76.200 57.430 76.220 ;
        RECT 58.400 76.200 59.100 76.400 ;
        RECT 69.200 76.200 69.400 81.900 ;
        RECT 57.200 75.700 58.000 76.200 ;
        RECT 57.200 75.680 57.430 75.700 ;
        RECT 49.040 75.300 57.040 75.420 ;
        RECT 48.000 75.190 57.040 75.300 ;
        RECT 48.000 75.100 49.300 75.190 ;
        RECT 48.000 70.500 48.200 75.100 ;
        RECT 48.400 74.300 48.900 74.800 ;
        RECT 58.400 74.300 58.600 76.200 ;
        RECT 65.400 76.150 69.400 76.200 ;
        RECT 60.975 76.000 69.400 76.150 ;
        RECT 60.975 75.920 65.665 76.000 ;
        RECT 69.200 75.600 69.400 76.000 ;
        RECT 66.800 75.580 69.400 75.600 ;
        RECT 59.140 75.400 69.400 75.580 ;
        RECT 59.140 75.350 67.140 75.400 ;
        RECT 67.400 75.090 68.300 75.100 ;
        RECT 67.345 74.600 68.300 75.090 ;
        RECT 67.345 74.550 67.575 74.600 ;
        RECT 48.400 73.920 48.600 74.300 ;
        RECT 56.800 74.280 58.600 74.300 ;
        RECT 49.040 74.100 58.600 74.280 ;
        RECT 49.040 74.050 57.040 74.100 ;
        RECT 48.400 73.120 48.680 73.920 ;
        RECT 57.800 73.800 58.000 74.100 ;
        RECT 59.140 74.060 67.140 74.290 ;
        RECT 57.300 73.790 58.000 73.800 ;
        RECT 57.200 73.300 58.000 73.790 ;
        RECT 57.200 73.250 57.430 73.300 ;
        RECT 59.200 73.150 59.400 74.060 ;
        RECT 60.980 73.700 65.670 73.720 ;
        RECT 69.200 73.700 69.400 75.400 ;
        RECT 60.980 73.500 69.400 73.700 ;
        RECT 60.980 73.490 65.670 73.500 ;
        RECT 48.400 72.900 48.600 73.120 ;
        RECT 49.040 72.900 57.040 72.990 ;
        RECT 59.145 72.920 67.145 73.150 ;
        RECT 48.400 72.760 57.040 72.900 ;
        RECT 48.400 72.700 49.300 72.760 ;
        RECT 67.400 72.660 68.300 72.700 ;
        RECT 48.400 71.800 48.900 72.300 ;
        RECT 67.350 72.200 68.300 72.660 ;
        RECT 58.200 71.900 58.700 72.200 ;
        RECT 67.350 72.120 67.600 72.200 ;
        RECT 56.800 71.850 58.700 71.900 ;
        RECT 48.400 71.490 48.600 71.800 ;
        RECT 49.040 71.700 58.700 71.850 ;
        RECT 49.040 71.620 57.040 71.700 ;
        RECT 48.400 71.300 48.680 71.490 ;
        RECT 48.450 70.690 48.680 71.300 ;
        RECT 57.200 71.300 57.430 71.360 ;
        RECT 57.200 70.820 58.000 71.300 ;
        RECT 57.300 70.800 58.000 70.820 ;
        RECT 49.040 70.500 57.040 70.560 ;
        RECT 48.000 70.330 57.040 70.500 ;
        RECT 48.000 70.300 49.300 70.330 ;
        RECT 48.000 68.100 48.200 70.300 ;
        RECT 48.400 69.400 48.900 69.900 ;
        RECT 58.200 69.500 58.400 71.700 ;
        RECT 59.145 71.630 67.145 71.860 ;
        RECT 59.200 70.170 59.400 71.630 ;
        RECT 60.975 70.510 65.645 70.740 ;
        RECT 67.400 70.200 67.600 72.120 ;
        RECT 66.900 70.170 67.600 70.200 ;
        RECT 59.155 70.000 67.600 70.170 ;
        RECT 59.155 69.940 67.155 70.000 ;
        RECT 68.500 69.700 69.000 69.900 ;
        RECT 67.400 69.680 69.000 69.700 ;
        RECT 56.800 69.420 58.400 69.500 ;
        RECT 48.400 69.060 48.600 69.400 ;
        RECT 49.040 69.300 58.400 69.420 ;
        RECT 49.040 69.190 57.040 69.300 ;
        RECT 48.400 68.900 48.680 69.060 ;
        RECT 48.450 68.260 48.680 68.900 ;
        RECT 57.200 68.900 57.430 68.930 ;
        RECT 57.200 68.400 58.000 68.900 ;
        RECT 58.200 68.800 58.400 69.300 ;
        RECT 67.315 69.400 69.000 69.680 ;
        RECT 67.315 69.140 67.545 69.400 ;
        RECT 59.155 68.800 67.155 68.880 ;
        RECT 58.200 68.650 67.155 68.800 ;
        RECT 58.200 68.600 59.400 68.650 ;
        RECT 57.200 68.390 57.430 68.400 ;
        RECT 49.040 68.100 57.040 68.130 ;
        RECT 48.000 67.900 57.040 68.100 ;
        RECT 48.000 65.600 48.200 67.900 ;
        RECT 48.400 66.900 48.900 67.400 ;
        RECT 58.200 67.000 58.400 68.600 ;
        RECT 69.200 67.800 69.400 73.500 ;
        RECT 65.400 67.750 69.400 67.800 ;
        RECT 60.975 67.600 69.400 67.750 ;
        RECT 60.975 67.520 65.665 67.600 ;
        RECT 69.200 67.200 69.400 67.600 ;
        RECT 66.800 67.180 69.400 67.200 ;
        RECT 56.800 66.990 58.400 67.000 ;
        RECT 48.400 66.630 48.600 66.900 ;
        RECT 49.040 66.800 58.400 66.990 ;
        RECT 59.140 67.000 69.400 67.180 ;
        RECT 59.140 66.950 67.140 67.000 ;
        RECT 49.040 66.760 57.040 66.800 ;
        RECT 48.400 66.400 48.680 66.630 ;
        RECT 48.450 65.830 48.680 66.400 ;
        RECT 57.200 66.000 58.000 66.500 ;
        RECT 57.200 65.960 57.430 66.000 ;
        RECT 49.040 65.600 57.040 65.700 ;
        RECT 48.000 65.470 57.040 65.600 ;
        RECT 48.000 65.400 49.300 65.470 ;
        RECT 48.000 63.200 48.200 65.400 ;
        RECT 48.400 64.500 48.900 65.000 ;
        RECT 58.200 64.600 58.400 66.800 ;
        RECT 67.400 66.690 68.300 66.700 ;
        RECT 67.345 66.200 68.300 66.690 ;
        RECT 67.345 66.150 67.575 66.200 ;
        RECT 59.140 65.660 67.140 65.890 ;
        RECT 59.300 64.780 59.500 65.660 ;
        RECT 69.200 65.400 69.400 67.000 ;
        RECT 65.400 65.350 69.400 65.400 ;
        RECT 60.975 65.200 69.400 65.350 ;
        RECT 60.975 65.120 65.665 65.200 ;
        RECT 56.800 64.560 58.400 64.600 ;
        RECT 48.400 64.200 48.600 64.500 ;
        RECT 49.040 64.400 58.400 64.560 ;
        RECT 59.140 64.550 67.140 64.780 ;
        RECT 49.040 64.330 57.040 64.400 ;
        RECT 67.400 64.290 68.300 64.300 ;
        RECT 48.400 63.900 48.680 64.200 ;
        RECT 57.300 64.070 58.000 64.100 ;
        RECT 48.450 63.400 48.680 63.900 ;
        RECT 57.200 63.600 58.000 64.070 ;
        RECT 67.345 63.800 68.300 64.290 ;
        RECT 67.345 63.750 67.575 63.800 ;
        RECT 57.200 63.530 57.430 63.600 ;
        RECT 59.140 63.400 67.140 63.490 ;
        RECT 49.040 63.200 57.040 63.270 ;
        RECT 48.000 63.040 57.040 63.200 ;
        RECT 58.200 63.260 67.140 63.400 ;
        RECT 58.200 63.200 59.400 63.260 ;
        RECT 48.000 63.000 49.300 63.040 ;
        RECT 48.000 53.700 48.200 63.000 ;
        RECT 48.400 62.500 53.200 62.700 ;
        RECT 48.400 62.100 48.900 62.500 ;
        RECT 50.700 62.100 50.900 62.500 ;
        RECT 48.400 62.080 49.400 62.100 ;
        RECT 50.700 62.080 51.700 62.100 ;
        RECT 48.400 61.900 50.040 62.080 ;
        RECT 48.400 60.195 48.600 61.900 ;
        RECT 49.040 61.850 50.040 61.900 ;
        RECT 50.700 61.900 52.340 62.080 ;
        RECT 50.700 60.195 50.900 61.900 ;
        RECT 51.340 61.850 52.340 61.900 ;
        RECT 53.000 60.195 53.200 62.500 ;
        RECT 54.300 62.080 56.200 62.100 ;
        RECT 53.640 61.900 56.940 62.080 ;
        RECT 53.640 61.850 54.640 61.900 ;
        RECT 55.940 61.850 56.940 61.900 ;
        RECT 48.400 59.900 48.680 60.195 ;
        RECT 50.700 59.900 50.980 60.195 ;
        RECT 53.000 59.900 53.280 60.195 ;
        RECT 48.450 55.445 48.680 59.900 ;
        RECT 50.200 55.800 50.430 59.840 ;
        RECT 49.040 53.700 50.040 53.790 ;
        RECT 48.000 53.560 50.040 53.700 ;
        RECT 48.000 53.500 49.300 53.560 ;
        RECT 49.000 53.300 49.300 53.500 ;
        RECT 49.000 52.800 49.500 53.300 ;
        RECT 50.200 52.600 50.400 55.800 ;
        RECT 50.750 55.445 50.980 59.900 ;
        RECT 52.500 55.800 52.730 59.840 ;
        RECT 51.340 53.560 52.340 53.790 ;
        RECT 51.400 53.300 51.700 53.560 ;
        RECT 51.400 52.800 51.900 53.300 ;
        RECT 52.500 52.600 52.700 55.800 ;
        RECT 53.050 55.700 53.280 59.900 ;
        RECT 54.800 55.800 55.030 59.840 ;
        RECT 53.050 55.445 53.300 55.700 ;
        RECT 53.100 53.300 53.300 55.445 ;
        RECT 53.640 53.560 54.640 53.790 ;
        RECT 53.700 53.300 54.000 53.560 ;
        RECT 53.100 53.100 53.500 53.300 ;
        RECT 50.200 52.100 50.700 52.600 ;
        RECT 52.500 52.100 53.000 52.600 ;
        RECT 53.300 51.900 53.500 53.100 ;
        RECT 53.700 52.800 54.200 53.300 ;
        RECT 54.800 52.600 55.000 55.800 ;
        RECT 54.700 52.100 55.200 52.600 ;
        RECT 55.350 51.900 55.580 58.920 ;
        RECT 53.300 51.700 55.580 51.900 ;
        RECT 35.740 50.720 44.100 50.800 ;
        RECT 39.400 50.600 44.100 50.720 ;
        RECT 38.020 48.500 38.520 49.000 ;
        RECT 38.020 48.250 38.220 48.500 ;
        RECT 35.980 48.020 40.020 48.250 ;
        RECT 33.720 47.600 33.970 47.860 ;
        RECT 42.030 47.700 42.260 47.860 ;
        RECT 33.740 47.440 33.970 47.600 ;
        RECT 42.020 47.440 42.260 47.700 ;
        RECT 33.120 46.900 33.320 47.365 ;
        RECT 42.020 46.900 42.220 47.440 ;
        RECT 33.120 46.700 43.720 46.900 ;
        RECT 39.220 45.995 43.320 46.000 ;
        RECT 32.620 45.500 32.900 45.980 ;
        RECT 35.480 45.800 43.320 45.995 ;
        RECT 35.480 45.765 39.520 45.800 ;
        RECT 33.240 45.500 33.470 45.560 ;
        RECT 32.620 45.300 33.470 45.500 ;
        RECT 41.530 45.400 41.760 45.560 ;
        RECT 32.670 45.080 32.900 45.300 ;
        RECT 33.240 45.140 33.470 45.300 ;
        RECT 41.520 45.200 42.920 45.400 ;
        RECT 41.530 45.140 41.760 45.200 ;
        RECT 42.720 44.000 42.920 45.200 ;
        RECT 42.420 43.700 42.920 44.000 ;
        RECT 41.420 43.640 42.920 43.700 ;
        RECT 33.760 43.500 42.920 43.640 ;
        RECT 33.760 43.410 41.760 43.500 ;
        RECT 33.170 42.800 33.400 43.280 ;
        RECT 41.920 43.100 42.150 43.150 ;
        RECT 43.120 43.100 43.320 45.800 ;
        RECT 41.920 42.900 43.320 43.100 ;
        RECT 33.170 42.480 33.420 42.800 ;
        RECT 41.920 42.610 42.150 42.900 ;
        RECT 42.420 42.600 42.920 42.900 ;
        RECT 27.320 41.400 27.520 42.140 ;
        RECT 33.220 41.800 33.420 42.480 ;
        RECT 33.760 42.120 41.760 42.350 ;
        RECT 33.820 41.800 34.020 42.120 ;
        RECT 43.520 41.800 43.720 46.700 ;
        RECT 33.220 41.600 43.720 41.800 ;
        RECT 43.900 46.800 44.100 50.600 ;
        RECT 54.600 47.500 54.800 51.700 ;
        RECT 55.350 51.620 55.580 51.700 ;
        RECT 57.100 51.975 57.330 58.565 ;
        RECT 57.100 48.700 57.300 51.975 ;
        RECT 58.200 48.700 58.400 63.200 ;
        RECT 69.200 63.000 69.400 65.200 ;
        RECT 65.400 62.950 69.400 63.000 ;
        RECT 60.975 62.800 69.400 62.950 ;
        RECT 60.975 62.720 65.665 62.800 ;
        RECT 69.200 62.400 69.400 62.800 ;
        RECT 66.800 62.380 69.400 62.400 ;
        RECT 59.140 62.200 69.400 62.380 ;
        RECT 59.140 62.150 67.140 62.200 ;
        RECT 67.400 61.890 68.300 61.900 ;
        RECT 67.345 61.400 68.300 61.890 ;
        RECT 67.345 61.350 67.575 61.400 ;
        RECT 59.140 60.860 67.140 61.090 ;
        RECT 59.200 59.985 59.400 60.860 ;
        RECT 69.200 60.600 69.400 62.200 ;
        RECT 65.400 60.555 69.400 60.600 ;
        RECT 60.975 60.400 69.400 60.555 ;
        RECT 60.975 60.325 65.665 60.400 ;
        RECT 59.140 59.755 67.140 59.985 ;
        RECT 67.400 59.495 68.300 59.500 ;
        RECT 67.345 59.000 68.300 59.495 ;
        RECT 67.345 58.955 67.575 59.000 ;
        RECT 59.140 58.600 67.140 58.695 ;
        RECT 68.500 58.600 69.000 58.800 ;
        RECT 59.140 58.465 69.000 58.600 ;
        RECT 66.900 58.400 69.000 58.465 ;
        RECT 68.500 58.300 69.000 58.400 ;
        RECT 69.200 58.100 69.400 60.400 ;
        RECT 62.300 58.050 69.400 58.100 ;
        RECT 62.080 57.900 69.400 58.050 ;
        RECT 62.080 57.820 62.980 57.900 ;
        RECT 59.480 57.500 60.280 57.550 ;
        RECT 56.600 48.690 58.400 48.700 ;
        RECT 55.940 48.500 58.400 48.690 ;
        RECT 58.600 57.320 60.280 57.500 ;
        RECT 62.300 57.480 62.500 57.820 ;
        RECT 63.700 57.550 64.700 57.600 ;
        RECT 58.600 57.300 59.800 57.320 ;
        RECT 58.600 56.900 58.800 57.300 ;
        RECT 62.140 57.250 62.560 57.480 ;
        RECT 63.700 57.400 65.245 57.550 ;
        RECT 59.120 56.900 59.350 56.960 ;
        RECT 58.600 56.700 59.350 56.900 ;
        RECT 55.940 48.460 56.940 48.500 ;
        RECT 56.000 48.200 56.200 48.460 ;
        RECT 56.000 47.700 56.500 48.200 ;
        RECT 58.600 47.500 58.800 56.700 ;
        RECT 59.120 48.960 59.350 56.700 ;
        RECT 60.410 49.300 60.640 56.960 ;
        RECT 62.765 51.500 62.995 55.240 ;
        RECT 62.765 51.200 63.000 51.500 ;
        RECT 60.410 48.960 60.700 49.300 ;
        RECT 62.200 49.190 62.400 49.200 ;
        RECT 62.140 48.960 62.560 49.190 ;
        RECT 59.610 48.570 60.150 48.800 ;
        RECT 59.900 48.300 60.100 48.570 ;
        RECT 59.600 47.800 60.100 48.300 ;
        RECT 60.500 48.300 60.700 48.960 ;
        RECT 60.500 48.000 61.000 48.300 ;
        RECT 62.200 48.000 62.400 48.960 ;
        RECT 60.500 47.800 62.400 48.000 ;
        RECT 54.600 47.300 58.800 47.500 ;
        RECT 59.900 47.600 60.100 47.800 ;
        RECT 62.800 47.600 63.000 51.200 ;
        RECT 59.900 47.400 63.000 47.600 ;
        RECT 63.700 48.700 63.900 57.400 ;
        RECT 64.365 57.320 65.245 57.400 ;
        RECT 67.800 57.000 68.300 57.300 ;
        RECT 64.600 56.980 68.300 57.000 ;
        RECT 64.440 56.800 68.300 56.980 ;
        RECT 68.500 56.800 69.000 57.300 ;
        RECT 64.440 56.750 64.860 56.800 ;
        RECT 68.600 55.100 68.800 56.800 ;
        RECT 65.020 52.700 65.250 54.740 ;
        RECT 65.020 52.500 66.000 52.700 ;
        RECT 65.020 50.700 65.250 52.500 ;
        RECT 65.500 52.200 66.000 52.500 ;
        RECT 67.720 51.400 67.950 55.100 ;
        RECT 67.600 51.100 67.950 51.400 ;
        RECT 68.510 54.800 68.800 55.100 ;
        RECT 68.510 51.100 68.740 54.800 ;
        RECT 69.200 54.265 69.400 57.900 ;
        RECT 69.080 53.900 69.400 54.265 ;
        RECT 69.080 51.575 69.310 53.900 ;
        RECT 63.700 48.690 64.700 48.700 ;
        RECT 63.700 48.500 64.860 48.690 ;
        RECT 58.600 47.200 58.800 47.300 ;
        RECT 63.700 47.200 63.900 48.500 ;
        RECT 64.440 48.460 64.860 48.500 ;
        RECT 58.600 47.000 63.900 47.200 ;
        RECT 67.600 46.800 67.800 51.100 ;
        RECT 68.000 50.665 68.460 50.895 ;
        RECT 68.100 49.900 68.300 50.665 ;
        RECT 68.100 49.200 68.800 49.900 ;
        RECT 68.100 48.200 68.800 48.900 ;
        RECT 43.900 46.600 67.800 46.800 ;
        RECT 18.520 41.200 26.320 41.400 ;
        RECT 27.320 41.200 42.220 41.400 ;
        RECT 14.520 40.430 15.020 41.000 ;
        RECT 16.420 40.800 17.420 41.000 ;
        RECT 14.500 40.200 15.040 40.430 ;
        RECT 16.420 40.040 16.620 40.800 ;
        RECT 16.920 40.430 17.420 40.800 ;
        RECT 16.920 40.300 17.470 40.430 ;
        RECT 16.930 40.200 17.470 40.300 ;
        RECT 18.820 40.040 19.020 41.200 ;
        RECT 19.420 40.430 19.920 41.000 ;
        RECT 19.360 40.300 19.920 40.430 ;
        RECT 19.360 40.200 19.900 40.300 ;
        RECT 21.220 40.040 21.420 41.200 ;
        RECT 21.820 40.430 22.320 41.000 ;
        RECT 21.790 40.200 22.330 40.430 ;
        RECT 23.720 40.040 23.920 41.200 ;
        RECT 24.220 40.430 24.720 41.000 ;
        RECT 24.220 40.200 24.760 40.430 ;
        RECT 26.120 40.040 26.320 41.200 ;
        RECT 26.620 40.430 27.120 41.000 ;
        RECT 26.620 40.300 27.190 40.430 ;
        RECT 26.650 40.200 27.190 40.300 ;
        RECT 32.155 40.300 38.745 40.330 ;
        RECT 42.020 40.300 42.220 41.200 ;
        RECT 32.155 40.100 42.220 40.300 ;
        RECT 6.620 39.800 6.950 40.040 ;
        RECT 6.720 32.040 6.950 39.800 ;
        RECT 8.010 32.300 8.240 40.040 ;
        RECT 9.120 39.800 9.380 40.040 ;
        RECT 8.010 32.040 8.320 32.300 ;
        RECT 9.150 32.040 9.380 39.800 ;
        RECT 10.440 32.300 10.670 40.040 ;
        RECT 11.520 39.800 11.810 40.040 ;
        RECT 10.440 32.040 10.720 32.300 ;
        RECT 11.580 32.040 11.810 39.800 ;
        RECT 12.870 32.300 13.100 40.040 ;
        RECT 13.920 39.800 14.240 40.040 ;
        RECT 12.870 32.040 13.120 32.300 ;
        RECT 14.010 32.040 14.240 39.800 ;
        RECT 15.300 32.300 15.530 40.040 ;
        RECT 16.420 39.800 16.670 40.040 ;
        RECT 15.300 32.040 15.620 32.300 ;
        RECT 16.440 32.040 16.670 39.800 ;
        RECT 17.730 32.300 17.960 40.040 ;
        RECT 18.820 39.800 19.100 40.040 ;
        RECT 17.730 32.040 18.020 32.300 ;
        RECT 18.870 32.040 19.100 39.800 ;
        RECT 20.160 32.300 20.390 40.040 ;
        RECT 21.220 39.800 21.530 40.040 ;
        RECT 20.160 32.040 20.420 32.300 ;
        RECT 21.300 32.040 21.530 39.800 ;
        RECT 22.590 32.040 22.820 40.040 ;
        RECT 23.720 39.800 23.960 40.040 ;
        RECT 23.730 32.040 23.960 39.800 ;
        RECT 25.020 32.300 25.250 40.040 ;
        RECT 26.120 39.800 26.390 40.040 ;
        RECT 25.020 32.040 25.320 32.300 ;
        RECT 26.160 32.040 26.390 39.800 ;
        RECT 27.450 32.300 27.680 40.040 ;
        RECT 42.020 39.940 42.220 40.100 ;
        RECT 28.640 39.200 28.870 39.940 ;
        RECT 42.020 39.600 42.260 39.940 ;
        RECT 28.620 38.940 28.870 39.200 ;
        RECT 42.030 39.200 42.260 39.600 ;
        RECT 42.520 39.200 43.020 39.500 ;
        RECT 42.030 39.000 43.020 39.200 ;
        RECT 42.030 38.940 42.260 39.000 ;
        RECT 28.620 37.640 28.820 38.940 ;
        RECT 31.800 38.350 39.100 38.580 ;
        RECT 30.880 38.000 34.920 38.030 ;
        RECT 38.120 38.000 38.620 38.200 ;
        RECT 30.880 37.800 38.620 38.000 ;
        RECT 38.120 37.700 38.620 37.800 ;
        RECT 38.820 37.800 39.020 38.350 ;
        RECT 43.220 37.800 43.420 41.600 ;
        RECT 28.620 37.300 28.870 37.640 ;
        RECT 28.640 36.640 28.870 37.300 ;
        RECT 36.930 37.000 37.160 37.640 ;
        RECT 38.820 37.600 43.420 37.800 ;
        RECT 37.420 37.000 37.920 37.200 ;
        RECT 36.930 36.700 37.920 37.000 ;
        RECT 36.930 36.640 37.160 36.700 ;
        RECT 38.820 36.500 39.020 37.600 ;
        RECT 37.420 36.300 39.020 36.500 ;
        RECT 35.020 36.280 37.620 36.300 ;
        RECT 30.525 36.200 37.620 36.280 ;
        RECT 28.020 36.100 37.620 36.200 ;
        RECT 28.020 36.050 35.275 36.100 ;
        RECT 28.020 36.000 30.820 36.050 ;
        RECT 28.020 33.900 28.220 36.000 ;
        RECT 30.880 35.700 34.920 35.730 ;
        RECT 38.120 35.700 38.620 36.000 ;
        RECT 30.880 35.500 38.620 35.700 ;
        RECT 28.640 34.700 28.870 35.340 ;
        RECT 28.620 34.340 28.870 34.700 ;
        RECT 36.930 34.700 37.160 35.340 ;
        RECT 37.420 34.700 37.920 34.900 ;
        RECT 36.930 34.400 37.920 34.700 ;
        RECT 36.930 34.340 37.160 34.400 ;
        RECT 28.620 33.900 28.820 34.340 ;
        RECT 30.525 33.900 35.275 33.980 ;
        RECT 28.020 33.750 35.275 33.900 ;
        RECT 28.020 33.700 30.820 33.750 ;
        RECT 27.450 32.040 27.720 32.300 ;
        RECT 6.220 31.600 6.720 31.900 ;
        RECT 7.080 31.600 7.880 31.680 ;
        RECT 6.220 31.450 7.880 31.600 ;
        RECT 6.220 31.400 7.220 31.450 ;
        RECT 8.120 31.200 8.320 32.040 ;
        RECT 8.720 31.600 9.220 31.900 ;
        RECT 9.510 31.600 10.310 31.680 ;
        RECT 8.720 31.450 10.310 31.600 ;
        RECT 8.720 31.400 9.720 31.450 ;
        RECT 10.520 31.200 10.720 32.040 ;
        RECT 11.120 31.600 11.620 31.900 ;
        RECT 11.940 31.600 12.740 31.680 ;
        RECT 11.120 31.450 12.740 31.600 ;
        RECT 11.120 31.400 12.120 31.450 ;
        RECT 12.920 31.200 13.120 32.040 ;
        RECT 13.520 31.600 14.020 31.900 ;
        RECT 14.370 31.600 15.170 31.680 ;
        RECT 13.520 31.450 15.170 31.600 ;
        RECT 13.520 31.400 14.620 31.450 ;
        RECT 15.420 31.200 15.620 32.040 ;
        RECT 15.920 31.600 16.420 31.900 ;
        RECT 16.800 31.600 17.600 31.680 ;
        RECT 17.820 31.600 18.020 32.040 ;
        RECT 15.920 31.400 18.020 31.600 ;
        RECT 18.420 31.600 18.920 31.900 ;
        RECT 19.230 31.600 20.030 31.680 ;
        RECT 18.420 31.450 20.030 31.600 ;
        RECT 18.420 31.400 19.420 31.450 ;
        RECT 20.220 31.200 20.420 32.040 ;
        RECT 20.820 31.600 21.320 31.900 ;
        RECT 21.660 31.600 22.460 31.680 ;
        RECT 20.820 31.450 22.460 31.600 ;
        RECT 20.820 31.400 21.820 31.450 ;
        RECT 22.620 31.200 22.820 32.040 ;
        RECT 23.320 31.600 23.820 31.900 ;
        RECT 24.090 31.600 24.890 31.680 ;
        RECT 23.320 31.450 24.890 31.600 ;
        RECT 23.320 31.400 24.320 31.450 ;
        RECT 25.120 31.200 25.320 32.040 ;
        RECT 25.720 31.600 26.220 31.900 ;
        RECT 26.520 31.600 27.320 31.680 ;
        RECT 25.720 31.450 27.320 31.600 ;
        RECT 25.720 31.400 26.820 31.450 ;
        RECT 27.520 31.200 27.720 32.040 ;
        RECT 28.020 31.900 28.220 33.700 ;
        RECT 30.880 33.400 34.920 33.430 ;
        RECT 38.120 33.400 38.620 33.700 ;
        RECT 30.880 33.200 38.620 33.400 ;
        RECT 28.640 32.400 28.870 33.040 ;
        RECT 28.620 32.040 28.870 32.400 ;
        RECT 36.930 32.300 37.160 33.040 ;
        RECT 37.420 32.300 37.920 32.500 ;
        RECT 36.930 32.040 37.920 32.300 ;
        RECT 28.620 31.900 28.820 32.040 ;
        RECT 28.020 31.600 28.820 31.900 ;
        RECT 37.020 32.000 37.920 32.040 ;
        RECT 30.525 31.600 35.275 31.680 ;
        RECT 28.020 31.450 35.275 31.600 ;
        RECT 28.020 31.400 30.820 31.450 ;
        RECT 37.020 31.200 37.220 32.000 ;
        RECT 8.120 31.000 37.220 31.200 ;
        RECT 2.300 26.310 36.900 26.400 ;
        RECT 2.300 26.200 39.265 26.310 ;
        RECT 2.300 25.700 3.000 26.200 ;
        RECT 6.220 22.665 6.420 26.200 ;
        RECT 6.720 24.140 6.920 26.200 ;
        RECT 7.220 24.575 7.720 25.300 ;
        RECT 7.220 24.400 7.770 24.575 ;
        RECT 7.230 24.345 7.770 24.400 ;
        RECT 6.720 23.800 6.970 24.140 ;
        RECT 6.170 22.400 6.420 22.665 ;
        RECT 6.170 17.975 6.400 22.400 ;
        RECT 6.740 16.140 6.970 23.800 ;
        RECT 8.030 16.400 8.260 24.140 ;
        RECT 8.620 22.665 8.820 26.200 ;
        RECT 12.120 25.500 12.620 26.000 ;
        RECT 9.720 24.575 10.220 25.300 ;
        RECT 9.660 24.400 10.220 24.575 ;
        RECT 12.120 24.600 12.320 25.500 ;
        RECT 12.120 24.530 12.820 24.600 ;
        RECT 12.120 24.400 13.170 24.530 ;
        RECT 9.660 24.345 10.200 24.400 ;
        RECT 12.120 24.140 12.320 24.400 ;
        RECT 12.630 24.300 13.170 24.400 ;
        RECT 8.600 17.975 8.830 22.665 ;
        RECT 9.170 16.400 9.400 24.140 ;
        RECT 8.030 16.200 9.400 16.400 ;
        RECT 8.030 16.140 8.260 16.200 ;
        RECT 9.170 16.140 9.400 16.200 ;
        RECT 10.460 16.400 10.690 24.140 ;
        RECT 12.120 23.900 12.370 24.140 ;
        RECT 11.570 22.600 11.800 22.630 ;
        RECT 11.570 22.400 11.820 22.600 ;
        RECT 11.570 17.960 11.800 22.400 ;
        RECT 12.140 16.400 12.370 23.900 ;
        RECT 10.460 16.200 12.370 16.400 ;
        RECT 10.460 16.140 10.690 16.200 ;
        RECT 12.140 16.140 12.370 16.200 ;
        RECT 13.430 16.400 13.660 24.140 ;
        RECT 14.520 22.665 14.720 26.200 ;
        RECT 15.120 24.140 15.320 26.200 ;
        RECT 15.620 24.575 16.120 25.300 ;
        RECT 15.620 24.400 16.170 24.575 ;
        RECT 15.630 24.345 16.170 24.400 ;
        RECT 15.120 23.800 15.370 24.140 ;
        RECT 14.520 22.400 14.800 22.665 ;
        RECT 14.570 17.975 14.800 22.400 ;
        RECT 13.430 16.140 13.720 16.400 ;
        RECT 15.140 16.140 15.370 23.800 ;
        RECT 16.430 16.400 16.660 24.140 ;
        RECT 17.020 22.670 17.220 26.200 ;
        RECT 20.820 25.500 21.320 26.000 ;
        RECT 18.020 24.600 18.520 25.300 ;
        RECT 18.020 24.400 20.720 24.600 ;
        RECT 21.020 24.545 21.320 25.500 ;
        RECT 21.020 24.400 21.580 24.545 ;
        RECT 18.060 24.350 18.600 24.400 ;
        RECT 20.520 24.155 20.720 24.400 ;
        RECT 21.040 24.315 21.580 24.400 ;
        RECT 17.000 17.980 17.230 22.670 ;
        RECT 17.570 16.400 17.800 24.145 ;
        RECT 16.430 16.200 17.800 16.400 ;
        RECT 16.430 16.140 16.660 16.200 ;
        RECT 17.570 16.145 17.800 16.200 ;
        RECT 18.860 16.400 19.090 24.145 ;
        RECT 20.520 23.900 20.780 24.155 ;
        RECT 19.980 17.975 20.210 22.645 ;
        RECT 20.550 16.400 20.780 23.900 ;
        RECT 18.860 16.200 20.780 16.400 ;
        RECT 18.860 16.145 19.090 16.200 ;
        RECT 20.550 16.155 20.780 16.200 ;
        RECT 21.840 16.400 22.070 24.155 ;
        RECT 22.920 22.665 23.120 26.200 ;
        RECT 23.520 24.140 23.720 26.200 ;
        RECT 24.020 24.575 24.520 25.300 ;
        RECT 24.020 24.400 24.570 24.575 ;
        RECT 24.030 24.345 24.570 24.400 ;
        RECT 23.520 23.800 23.770 24.140 ;
        RECT 22.920 22.400 23.200 22.665 ;
        RECT 22.970 17.975 23.200 22.400 ;
        RECT 21.840 16.155 22.120 16.400 ;
        RECT 13.520 16.100 13.720 16.140 ;
        RECT 13.520 15.900 14.520 16.100 ;
        RECT 13.620 15.400 14.120 15.700 ;
        RECT 14.320 15.600 14.520 15.900 ;
        RECT 14.320 15.400 16.620 15.600 ;
        RECT 6.620 15.200 14.120 15.400 ;
        RECT 6.620 14.040 6.820 15.200 ;
        RECT 7.220 14.430 7.720 15.000 ;
        RECT 7.210 14.200 7.750 14.430 ;
        RECT 9.120 14.040 9.320 15.200 ;
        RECT 9.620 14.430 10.120 15.000 ;
        RECT 9.620 14.300 10.180 14.430 ;
        RECT 9.640 14.200 10.180 14.300 ;
        RECT 11.520 14.040 11.720 15.200 ;
        RECT 12.020 14.430 12.520 15.000 ;
        RECT 12.020 14.300 12.610 14.430 ;
        RECT 12.070 14.200 12.610 14.300 ;
        RECT 13.920 14.040 14.120 15.200 ;
        RECT 16.420 15.000 16.620 15.400 ;
        RECT 18.520 15.400 19.020 15.700 ;
        RECT 21.920 15.400 22.120 16.155 ;
        RECT 23.540 16.140 23.770 23.800 ;
        RECT 24.830 16.500 25.060 24.140 ;
        RECT 25.320 22.665 25.520 26.200 ;
        RECT 26.420 24.575 26.920 25.300 ;
        RECT 26.420 24.400 26.970 24.575 ;
        RECT 26.430 24.345 26.970 24.400 ;
        RECT 25.320 22.400 25.600 22.665 ;
        RECT 25.370 17.975 25.600 22.400 ;
        RECT 25.940 16.500 26.170 24.140 ;
        RECT 24.830 16.300 26.170 16.500 ;
        RECT 24.830 16.140 25.060 16.300 ;
        RECT 25.940 16.140 26.170 16.300 ;
        RECT 27.230 16.400 27.460 24.140 ;
        RECT 27.720 22.665 27.920 26.200 ;
        RECT 28.320 24.140 28.520 26.200 ;
        RECT 28.820 24.575 29.320 25.300 ;
        RECT 28.820 24.400 29.370 24.575 ;
        RECT 28.830 24.345 29.370 24.400 ;
        RECT 28.320 23.800 28.570 24.140 ;
        RECT 27.720 22.400 28.000 22.665 ;
        RECT 27.770 17.975 28.000 22.400 ;
        RECT 27.230 16.140 27.520 16.400 ;
        RECT 28.340 16.140 28.570 23.800 ;
        RECT 29.630 16.400 29.860 24.140 ;
        RECT 30.120 22.665 30.320 26.200 ;
        RECT 32.600 26.100 32.820 26.200 ;
        RECT 35.000 26.100 39.265 26.200 ;
        RECT 31.920 25.500 32.420 26.000 ;
        RECT 31.220 24.575 31.720 25.300 ;
        RECT 31.220 24.400 31.765 24.575 ;
        RECT 31.225 24.345 31.765 24.400 ;
        RECT 32.120 24.140 32.320 25.500 ;
        RECT 30.120 22.400 30.395 22.665 ;
        RECT 30.165 17.975 30.395 22.400 ;
        RECT 30.735 16.400 30.965 24.140 ;
        RECT 29.630 16.200 30.965 16.400 ;
        RECT 29.630 16.140 29.860 16.200 ;
        RECT 30.735 16.140 30.965 16.200 ;
        RECT 32.025 23.900 32.320 24.140 ;
        RECT 32.025 16.140 32.255 23.900 ;
        RECT 32.620 19.980 32.820 26.100 ;
        RECT 36.575 26.080 39.265 26.100 ;
        RECT 33.400 25.800 33.900 26.000 ;
        RECT 33.400 25.740 36.000 25.800 ;
        RECT 33.400 25.600 39.740 25.740 ;
        RECT 33.400 25.500 33.900 25.600 ;
        RECT 35.740 25.510 39.740 25.600 ;
        RECT 39.945 25.300 40.175 25.460 ;
        RECT 40.900 25.300 41.600 25.800 ;
        RECT 33.420 24.800 33.920 25.300 ;
        RECT 39.945 25.100 41.600 25.300 ;
        RECT 41.900 25.100 42.600 25.800 ;
        RECT 39.945 25.000 40.175 25.100 ;
        RECT 33.170 21.700 33.400 22.245 ;
        RECT 33.120 21.365 33.400 21.700 ;
        RECT 33.720 21.860 33.920 24.800 ;
        RECT 35.740 24.900 39.740 24.950 ;
        RECT 35.740 24.800 39.800 24.900 ;
        RECT 43.900 24.800 44.100 46.600 ;
        RECT 60.975 42.500 65.665 42.550 ;
        RECT 71.000 42.500 73.000 84.300 ;
        RECT 48.400 42.000 48.900 42.500 ;
        RECT 60.975 42.320 73.000 42.500 ;
        RECT 65.400 42.300 73.000 42.320 ;
        RECT 56.800 42.000 58.400 42.100 ;
        RECT 69.200 42.000 69.400 42.300 ;
        RECT 48.400 41.640 48.600 42.000 ;
        RECT 49.040 41.900 58.400 42.000 ;
        RECT 66.800 41.980 69.400 42.000 ;
        RECT 49.040 41.770 57.040 41.900 ;
        RECT 48.400 41.500 48.680 41.640 ;
        RECT 48.450 40.840 48.680 41.500 ;
        RECT 57.200 41.500 57.430 41.510 ;
        RECT 57.200 41.000 58.000 41.500 ;
        RECT 57.200 40.970 57.430 41.000 ;
        RECT 49.040 40.600 57.040 40.710 ;
        RECT 35.740 24.720 44.100 24.800 ;
        RECT 39.400 24.600 44.100 24.720 ;
        RECT 38.020 22.500 38.520 23.000 ;
        RECT 38.020 22.250 38.220 22.500 ;
        RECT 35.980 22.020 40.020 22.250 ;
        RECT 33.720 21.600 33.970 21.860 ;
        RECT 42.030 21.700 42.260 21.860 ;
        RECT 33.740 21.440 33.970 21.600 ;
        RECT 42.020 21.440 42.260 21.700 ;
        RECT 33.120 20.900 33.320 21.365 ;
        RECT 42.020 20.900 42.220 21.440 ;
        RECT 33.120 20.700 43.720 20.900 ;
        RECT 39.220 19.995 43.320 20.000 ;
        RECT 32.620 19.500 32.900 19.980 ;
        RECT 35.480 19.800 43.320 19.995 ;
        RECT 35.480 19.765 39.520 19.800 ;
        RECT 33.240 19.500 33.470 19.560 ;
        RECT 32.620 19.300 33.470 19.500 ;
        RECT 41.530 19.400 41.760 19.560 ;
        RECT 32.670 19.080 32.900 19.300 ;
        RECT 33.240 19.140 33.470 19.300 ;
        RECT 41.520 19.200 42.920 19.400 ;
        RECT 41.530 19.140 41.760 19.200 ;
        RECT 42.720 18.000 42.920 19.200 ;
        RECT 42.420 17.700 42.920 18.000 ;
        RECT 41.420 17.640 42.920 17.700 ;
        RECT 33.760 17.500 42.920 17.640 ;
        RECT 33.760 17.410 41.760 17.500 ;
        RECT 33.170 16.800 33.400 17.280 ;
        RECT 41.920 17.100 42.150 17.150 ;
        RECT 43.120 17.100 43.320 19.800 ;
        RECT 41.920 16.900 43.320 17.100 ;
        RECT 33.170 16.480 33.420 16.800 ;
        RECT 41.920 16.610 42.150 16.900 ;
        RECT 42.420 16.600 42.920 16.900 ;
        RECT 27.320 15.400 27.520 16.140 ;
        RECT 33.220 15.800 33.420 16.480 ;
        RECT 33.760 16.120 41.760 16.350 ;
        RECT 33.820 15.800 34.020 16.120 ;
        RECT 43.520 15.800 43.720 20.700 ;
        RECT 33.220 15.600 43.720 15.800 ;
        RECT 18.520 15.200 26.320 15.400 ;
        RECT 27.320 15.200 42.220 15.400 ;
        RECT 14.520 14.430 15.020 15.000 ;
        RECT 16.420 14.800 17.420 15.000 ;
        RECT 14.500 14.200 15.040 14.430 ;
        RECT 16.420 14.040 16.620 14.800 ;
        RECT 16.920 14.430 17.420 14.800 ;
        RECT 16.920 14.300 17.470 14.430 ;
        RECT 16.930 14.200 17.470 14.300 ;
        RECT 18.820 14.040 19.020 15.200 ;
        RECT 19.420 14.430 19.920 15.000 ;
        RECT 19.360 14.300 19.920 14.430 ;
        RECT 19.360 14.200 19.900 14.300 ;
        RECT 21.220 14.040 21.420 15.200 ;
        RECT 21.820 14.430 22.320 15.000 ;
        RECT 21.790 14.200 22.330 14.430 ;
        RECT 23.720 14.040 23.920 15.200 ;
        RECT 24.220 14.430 24.720 15.000 ;
        RECT 24.220 14.200 24.760 14.430 ;
        RECT 26.120 14.040 26.320 15.200 ;
        RECT 26.620 14.430 27.120 15.000 ;
        RECT 26.620 14.300 27.190 14.430 ;
        RECT 26.650 14.200 27.190 14.300 ;
        RECT 32.155 14.300 38.745 14.330 ;
        RECT 42.020 14.300 42.220 15.200 ;
        RECT 32.155 14.100 42.220 14.300 ;
        RECT 6.620 13.800 6.950 14.040 ;
        RECT 6.720 6.040 6.950 13.800 ;
        RECT 8.010 6.300 8.240 14.040 ;
        RECT 9.120 13.800 9.380 14.040 ;
        RECT 8.010 6.040 8.320 6.300 ;
        RECT 9.150 6.040 9.380 13.800 ;
        RECT 10.440 6.300 10.670 14.040 ;
        RECT 11.520 13.800 11.810 14.040 ;
        RECT 10.440 6.040 10.720 6.300 ;
        RECT 11.580 6.040 11.810 13.800 ;
        RECT 12.870 6.300 13.100 14.040 ;
        RECT 13.920 13.800 14.240 14.040 ;
        RECT 12.870 6.040 13.120 6.300 ;
        RECT 14.010 6.040 14.240 13.800 ;
        RECT 15.300 6.300 15.530 14.040 ;
        RECT 16.420 13.800 16.670 14.040 ;
        RECT 15.300 6.040 15.620 6.300 ;
        RECT 16.440 6.040 16.670 13.800 ;
        RECT 17.730 6.300 17.960 14.040 ;
        RECT 18.820 13.800 19.100 14.040 ;
        RECT 17.730 6.040 18.020 6.300 ;
        RECT 18.870 6.040 19.100 13.800 ;
        RECT 20.160 6.300 20.390 14.040 ;
        RECT 21.220 13.800 21.530 14.040 ;
        RECT 20.160 6.040 20.420 6.300 ;
        RECT 21.300 6.040 21.530 13.800 ;
        RECT 22.590 6.040 22.820 14.040 ;
        RECT 23.720 13.800 23.960 14.040 ;
        RECT 23.730 6.040 23.960 13.800 ;
        RECT 25.020 6.300 25.250 14.040 ;
        RECT 26.120 13.800 26.390 14.040 ;
        RECT 25.020 6.040 25.320 6.300 ;
        RECT 26.160 6.040 26.390 13.800 ;
        RECT 27.450 6.300 27.680 14.040 ;
        RECT 42.020 13.940 42.220 14.100 ;
        RECT 28.640 13.200 28.870 13.940 ;
        RECT 42.020 13.600 42.260 13.940 ;
        RECT 28.620 12.940 28.870 13.200 ;
        RECT 42.030 13.200 42.260 13.600 ;
        RECT 42.520 13.200 43.020 13.500 ;
        RECT 42.030 13.000 43.020 13.200 ;
        RECT 42.030 12.940 42.260 13.000 ;
        RECT 28.620 11.640 28.820 12.940 ;
        RECT 31.800 12.350 39.100 12.580 ;
        RECT 30.880 12.000 34.920 12.030 ;
        RECT 38.120 12.000 38.620 12.200 ;
        RECT 30.880 11.800 38.620 12.000 ;
        RECT 38.120 11.700 38.620 11.800 ;
        RECT 38.820 11.800 39.020 12.350 ;
        RECT 43.220 11.800 43.420 15.600 ;
        RECT 28.620 11.300 28.870 11.640 ;
        RECT 28.640 10.640 28.870 11.300 ;
        RECT 36.930 11.000 37.160 11.640 ;
        RECT 38.820 11.600 43.420 11.800 ;
        RECT 37.420 11.000 37.920 11.200 ;
        RECT 36.930 10.700 37.920 11.000 ;
        RECT 36.930 10.640 37.160 10.700 ;
        RECT 38.820 10.500 39.020 11.600 ;
        RECT 37.420 10.300 39.020 10.500 ;
        RECT 35.020 10.280 37.620 10.300 ;
        RECT 30.525 10.200 37.620 10.280 ;
        RECT 28.020 10.100 37.620 10.200 ;
        RECT 28.020 10.050 35.275 10.100 ;
        RECT 28.020 10.000 30.820 10.050 ;
        RECT 28.020 7.900 28.220 10.000 ;
        RECT 30.880 9.700 34.920 9.730 ;
        RECT 38.120 9.700 38.620 10.000 ;
        RECT 30.880 9.500 38.620 9.700 ;
        RECT 28.640 8.700 28.870 9.340 ;
        RECT 28.620 8.340 28.870 8.700 ;
        RECT 36.930 8.700 37.160 9.340 ;
        RECT 37.420 8.700 37.920 8.900 ;
        RECT 36.930 8.400 37.920 8.700 ;
        RECT 36.930 8.340 37.160 8.400 ;
        RECT 28.620 7.900 28.820 8.340 ;
        RECT 30.525 7.900 35.275 7.980 ;
        RECT 28.020 7.750 35.275 7.900 ;
        RECT 28.020 7.700 30.820 7.750 ;
        RECT 27.450 6.040 27.720 6.300 ;
        RECT 6.220 5.600 6.720 5.900 ;
        RECT 7.080 5.600 7.880 5.680 ;
        RECT 6.220 5.450 7.880 5.600 ;
        RECT 6.220 5.400 7.220 5.450 ;
        RECT 8.120 5.200 8.320 6.040 ;
        RECT 8.720 5.600 9.220 5.900 ;
        RECT 9.510 5.600 10.310 5.680 ;
        RECT 8.720 5.450 10.310 5.600 ;
        RECT 8.720 5.400 9.720 5.450 ;
        RECT 10.520 5.200 10.720 6.040 ;
        RECT 11.120 5.600 11.620 5.900 ;
        RECT 11.940 5.600 12.740 5.680 ;
        RECT 11.120 5.450 12.740 5.600 ;
        RECT 11.120 5.400 12.120 5.450 ;
        RECT 12.920 5.200 13.120 6.040 ;
        RECT 13.520 5.600 14.020 5.900 ;
        RECT 14.370 5.600 15.170 5.680 ;
        RECT 13.520 5.450 15.170 5.600 ;
        RECT 13.520 5.400 14.620 5.450 ;
        RECT 15.420 5.200 15.620 6.040 ;
        RECT 15.920 5.600 16.420 5.900 ;
        RECT 16.800 5.600 17.600 5.680 ;
        RECT 17.820 5.600 18.020 6.040 ;
        RECT 15.920 5.400 18.020 5.600 ;
        RECT 18.420 5.600 18.920 5.900 ;
        RECT 19.230 5.600 20.030 5.680 ;
        RECT 18.420 5.450 20.030 5.600 ;
        RECT 18.420 5.400 19.420 5.450 ;
        RECT 20.220 5.200 20.420 6.040 ;
        RECT 20.820 5.600 21.320 5.900 ;
        RECT 21.660 5.600 22.460 5.680 ;
        RECT 20.820 5.450 22.460 5.600 ;
        RECT 20.820 5.400 21.820 5.450 ;
        RECT 22.620 5.200 22.820 6.040 ;
        RECT 23.320 5.600 23.820 5.900 ;
        RECT 24.090 5.600 24.890 5.680 ;
        RECT 23.320 5.450 24.890 5.600 ;
        RECT 23.320 5.400 24.320 5.450 ;
        RECT 25.120 5.200 25.320 6.040 ;
        RECT 25.720 5.600 26.220 5.900 ;
        RECT 26.520 5.600 27.320 5.680 ;
        RECT 25.720 5.450 27.320 5.600 ;
        RECT 25.720 5.400 26.820 5.450 ;
        RECT 27.520 5.200 27.720 6.040 ;
        RECT 28.020 5.900 28.220 7.700 ;
        RECT 30.880 7.400 34.920 7.430 ;
        RECT 38.120 7.400 38.620 7.700 ;
        RECT 30.880 7.200 38.620 7.400 ;
        RECT 28.640 6.400 28.870 7.040 ;
        RECT 28.620 6.040 28.870 6.400 ;
        RECT 36.930 6.300 37.160 7.040 ;
        RECT 37.420 6.300 37.920 6.500 ;
        RECT 36.930 6.040 37.920 6.300 ;
        RECT 28.620 5.900 28.820 6.040 ;
        RECT 28.020 5.600 28.820 5.900 ;
        RECT 37.020 6.000 37.920 6.040 ;
        RECT 30.525 5.600 35.275 5.680 ;
        RECT 28.020 5.450 35.275 5.600 ;
        RECT 28.020 5.400 30.820 5.450 ;
        RECT 37.020 5.200 37.220 6.000 ;
        RECT 8.120 5.000 37.220 5.200 ;
        RECT 43.900 4.800 44.100 24.600 ;
        RECT 48.000 40.480 57.040 40.600 ;
        RECT 48.000 40.400 49.300 40.480 ;
        RECT 48.000 38.200 48.200 40.400 ;
        RECT 48.400 39.500 48.900 40.000 ;
        RECT 58.200 39.600 58.400 41.900 ;
        RECT 59.140 41.800 69.400 41.980 ;
        RECT 59.140 41.750 67.140 41.800 ;
        RECT 67.400 41.490 68.300 41.500 ;
        RECT 67.345 41.000 68.300 41.490 ;
        RECT 67.345 40.950 67.575 41.000 ;
        RECT 59.140 40.460 67.140 40.690 ;
        RECT 56.800 39.570 58.400 39.600 ;
        RECT 48.400 39.210 48.600 39.500 ;
        RECT 49.040 39.400 58.400 39.570 ;
        RECT 59.200 39.550 59.400 40.460 ;
        RECT 60.975 40.100 65.665 40.120 ;
        RECT 69.200 40.100 69.400 41.800 ;
        RECT 60.975 39.900 69.400 40.100 ;
        RECT 60.975 39.890 65.665 39.900 ;
        RECT 49.040 39.340 57.040 39.400 ;
        RECT 48.400 39.000 48.680 39.210 ;
        RECT 57.300 39.080 58.000 39.100 ;
        RECT 48.450 38.410 48.680 39.000 ;
        RECT 57.200 38.600 58.000 39.080 ;
        RECT 57.200 38.540 57.430 38.600 ;
        RECT 49.040 38.200 57.040 38.280 ;
        RECT 48.000 38.050 57.040 38.200 ;
        RECT 48.000 38.000 49.300 38.050 ;
        RECT 48.000 35.800 48.200 38.000 ;
        RECT 48.400 37.100 48.900 37.600 ;
        RECT 58.200 37.200 58.400 39.400 ;
        RECT 59.140 39.320 67.140 39.550 ;
        RECT 67.345 39.000 67.575 39.060 ;
        RECT 67.345 38.520 68.300 39.000 ;
        RECT 67.400 38.500 68.300 38.520 ;
        RECT 59.140 38.030 67.140 38.260 ;
        RECT 56.800 37.140 58.400 37.200 ;
        RECT 48.400 36.780 48.600 37.100 ;
        RECT 49.040 37.000 58.400 37.140 ;
        RECT 49.040 36.910 57.040 37.000 ;
        RECT 48.400 36.600 48.680 36.780 ;
        RECT 57.300 36.650 58.000 36.700 ;
        RECT 48.450 35.980 48.680 36.600 ;
        RECT 57.200 36.200 58.000 36.650 ;
        RECT 57.200 36.110 57.430 36.200 ;
        RECT 49.040 35.800 57.040 35.850 ;
        RECT 48.000 35.620 57.040 35.800 ;
        RECT 48.000 35.600 49.300 35.620 ;
        RECT 48.000 33.300 48.200 35.600 ;
        RECT 48.400 34.700 48.900 35.200 ;
        RECT 58.200 35.100 58.400 37.000 ;
        RECT 59.200 36.580 59.400 38.030 ;
        RECT 60.960 36.920 65.630 37.150 ;
        RECT 65.400 36.900 65.600 36.920 ;
        RECT 66.900 36.580 69.000 36.600 ;
        RECT 59.140 36.400 69.000 36.580 ;
        RECT 59.140 36.350 67.140 36.400 ;
        RECT 67.400 36.090 67.600 36.400 ;
        RECT 68.500 36.100 69.000 36.400 ;
        RECT 67.300 35.900 67.600 36.090 ;
        RECT 67.300 35.550 67.530 35.900 ;
        RECT 59.140 35.200 67.140 35.290 ;
        RECT 58.200 34.800 58.700 35.100 ;
        RECT 56.800 34.710 58.700 34.800 ;
        RECT 48.400 34.350 48.600 34.700 ;
        RECT 49.040 34.600 58.700 34.710 ;
        RECT 58.900 35.060 67.140 35.200 ;
        RECT 58.900 35.000 59.400 35.060 ;
        RECT 49.040 34.480 57.040 34.600 ;
        RECT 58.900 34.400 59.100 35.000 ;
        RECT 48.400 34.100 48.680 34.350 ;
        RECT 48.450 33.550 48.680 34.100 ;
        RECT 57.200 34.200 57.430 34.220 ;
        RECT 58.400 34.200 59.100 34.400 ;
        RECT 69.200 34.200 69.400 39.900 ;
        RECT 57.200 33.700 58.000 34.200 ;
        RECT 57.200 33.680 57.430 33.700 ;
        RECT 49.040 33.300 57.040 33.420 ;
        RECT 48.000 33.190 57.040 33.300 ;
        RECT 48.000 33.100 49.300 33.190 ;
        RECT 48.000 28.500 48.200 33.100 ;
        RECT 48.400 32.300 48.900 32.800 ;
        RECT 58.400 32.300 58.600 34.200 ;
        RECT 65.400 34.150 69.400 34.200 ;
        RECT 60.975 34.000 69.400 34.150 ;
        RECT 60.975 33.920 65.665 34.000 ;
        RECT 69.200 33.600 69.400 34.000 ;
        RECT 66.800 33.580 69.400 33.600 ;
        RECT 59.140 33.400 69.400 33.580 ;
        RECT 59.140 33.350 67.140 33.400 ;
        RECT 67.400 33.090 68.300 33.100 ;
        RECT 67.345 32.600 68.300 33.090 ;
        RECT 67.345 32.550 67.575 32.600 ;
        RECT 48.400 31.920 48.600 32.300 ;
        RECT 56.800 32.280 58.600 32.300 ;
        RECT 49.040 32.100 58.600 32.280 ;
        RECT 49.040 32.050 57.040 32.100 ;
        RECT 48.400 31.120 48.680 31.920 ;
        RECT 57.800 31.800 58.000 32.100 ;
        RECT 59.140 32.060 67.140 32.290 ;
        RECT 57.300 31.790 58.000 31.800 ;
        RECT 57.200 31.300 58.000 31.790 ;
        RECT 57.200 31.250 57.430 31.300 ;
        RECT 59.200 31.150 59.400 32.060 ;
        RECT 60.980 31.700 65.670 31.720 ;
        RECT 69.200 31.700 69.400 33.400 ;
        RECT 60.980 31.500 69.400 31.700 ;
        RECT 60.980 31.490 65.670 31.500 ;
        RECT 48.400 30.900 48.600 31.120 ;
        RECT 49.040 30.900 57.040 30.990 ;
        RECT 59.145 30.920 67.145 31.150 ;
        RECT 48.400 30.760 57.040 30.900 ;
        RECT 48.400 30.700 49.300 30.760 ;
        RECT 67.400 30.660 68.300 30.700 ;
        RECT 48.400 29.800 48.900 30.300 ;
        RECT 67.350 30.200 68.300 30.660 ;
        RECT 58.200 29.900 58.700 30.200 ;
        RECT 67.350 30.120 67.600 30.200 ;
        RECT 56.800 29.850 58.700 29.900 ;
        RECT 48.400 29.490 48.600 29.800 ;
        RECT 49.040 29.700 58.700 29.850 ;
        RECT 49.040 29.620 57.040 29.700 ;
        RECT 48.400 29.300 48.680 29.490 ;
        RECT 48.450 28.690 48.680 29.300 ;
        RECT 57.200 29.300 57.430 29.360 ;
        RECT 57.200 28.820 58.000 29.300 ;
        RECT 57.300 28.800 58.000 28.820 ;
        RECT 49.040 28.500 57.040 28.560 ;
        RECT 48.000 28.330 57.040 28.500 ;
        RECT 48.000 28.300 49.300 28.330 ;
        RECT 48.000 26.100 48.200 28.300 ;
        RECT 48.400 27.400 48.900 27.900 ;
        RECT 58.200 27.500 58.400 29.700 ;
        RECT 59.145 29.630 67.145 29.860 ;
        RECT 59.200 28.170 59.400 29.630 ;
        RECT 60.975 28.510 65.645 28.740 ;
        RECT 67.400 28.200 67.600 30.120 ;
        RECT 66.900 28.170 67.600 28.200 ;
        RECT 59.155 28.000 67.600 28.170 ;
        RECT 59.155 27.940 67.155 28.000 ;
        RECT 68.500 27.700 69.000 27.900 ;
        RECT 67.400 27.680 69.000 27.700 ;
        RECT 56.800 27.420 58.400 27.500 ;
        RECT 48.400 27.060 48.600 27.400 ;
        RECT 49.040 27.300 58.400 27.420 ;
        RECT 49.040 27.190 57.040 27.300 ;
        RECT 48.400 26.900 48.680 27.060 ;
        RECT 48.450 26.260 48.680 26.900 ;
        RECT 57.200 26.900 57.430 26.930 ;
        RECT 57.200 26.400 58.000 26.900 ;
        RECT 58.200 26.800 58.400 27.300 ;
        RECT 67.315 27.400 69.000 27.680 ;
        RECT 67.315 27.140 67.545 27.400 ;
        RECT 59.155 26.800 67.155 26.880 ;
        RECT 58.200 26.650 67.155 26.800 ;
        RECT 58.200 26.600 59.400 26.650 ;
        RECT 57.200 26.390 57.430 26.400 ;
        RECT 49.040 26.100 57.040 26.130 ;
        RECT 48.000 25.900 57.040 26.100 ;
        RECT 48.000 23.600 48.200 25.900 ;
        RECT 48.400 24.900 48.900 25.400 ;
        RECT 58.200 25.000 58.400 26.600 ;
        RECT 69.200 25.800 69.400 31.500 ;
        RECT 65.400 25.750 69.400 25.800 ;
        RECT 60.975 25.600 69.400 25.750 ;
        RECT 60.975 25.520 65.665 25.600 ;
        RECT 69.200 25.200 69.400 25.600 ;
        RECT 66.800 25.180 69.400 25.200 ;
        RECT 56.800 24.990 58.400 25.000 ;
        RECT 48.400 24.630 48.600 24.900 ;
        RECT 49.040 24.800 58.400 24.990 ;
        RECT 59.140 25.000 69.400 25.180 ;
        RECT 59.140 24.950 67.140 25.000 ;
        RECT 49.040 24.760 57.040 24.800 ;
        RECT 48.400 24.400 48.680 24.630 ;
        RECT 48.450 23.830 48.680 24.400 ;
        RECT 57.200 24.000 58.000 24.500 ;
        RECT 57.200 23.960 57.430 24.000 ;
        RECT 49.040 23.600 57.040 23.700 ;
        RECT 48.000 23.470 57.040 23.600 ;
        RECT 48.000 23.400 49.300 23.470 ;
        RECT 48.000 21.200 48.200 23.400 ;
        RECT 48.400 22.500 48.900 23.000 ;
        RECT 58.200 22.600 58.400 24.800 ;
        RECT 67.400 24.690 68.300 24.700 ;
        RECT 67.345 24.200 68.300 24.690 ;
        RECT 67.345 24.150 67.575 24.200 ;
        RECT 59.140 23.660 67.140 23.890 ;
        RECT 59.300 22.780 59.500 23.660 ;
        RECT 69.200 23.400 69.400 25.000 ;
        RECT 65.400 23.350 69.400 23.400 ;
        RECT 60.975 23.200 69.400 23.350 ;
        RECT 60.975 23.120 65.665 23.200 ;
        RECT 56.800 22.560 58.400 22.600 ;
        RECT 48.400 22.200 48.600 22.500 ;
        RECT 49.040 22.400 58.400 22.560 ;
        RECT 59.140 22.550 67.140 22.780 ;
        RECT 49.040 22.330 57.040 22.400 ;
        RECT 67.400 22.290 68.300 22.300 ;
        RECT 48.400 21.900 48.680 22.200 ;
        RECT 57.300 22.070 58.000 22.100 ;
        RECT 48.450 21.400 48.680 21.900 ;
        RECT 57.200 21.600 58.000 22.070 ;
        RECT 67.345 21.800 68.300 22.290 ;
        RECT 67.345 21.750 67.575 21.800 ;
        RECT 57.200 21.530 57.430 21.600 ;
        RECT 59.140 21.400 67.140 21.490 ;
        RECT 49.040 21.200 57.040 21.270 ;
        RECT 48.000 21.040 57.040 21.200 ;
        RECT 58.200 21.260 67.140 21.400 ;
        RECT 58.200 21.200 59.400 21.260 ;
        RECT 48.000 21.000 49.300 21.040 ;
        RECT 48.000 11.700 48.200 21.000 ;
        RECT 48.400 20.500 53.200 20.700 ;
        RECT 48.400 20.100 48.900 20.500 ;
        RECT 50.700 20.100 50.900 20.500 ;
        RECT 48.400 20.080 49.400 20.100 ;
        RECT 50.700 20.080 51.700 20.100 ;
        RECT 48.400 19.900 50.040 20.080 ;
        RECT 48.400 18.195 48.600 19.900 ;
        RECT 49.040 19.850 50.040 19.900 ;
        RECT 50.700 19.900 52.340 20.080 ;
        RECT 50.700 18.195 50.900 19.900 ;
        RECT 51.340 19.850 52.340 19.900 ;
        RECT 53.000 18.195 53.200 20.500 ;
        RECT 54.300 20.080 56.200 20.100 ;
        RECT 53.640 19.900 56.940 20.080 ;
        RECT 53.640 19.850 54.640 19.900 ;
        RECT 55.940 19.850 56.940 19.900 ;
        RECT 48.400 17.900 48.680 18.195 ;
        RECT 50.700 17.900 50.980 18.195 ;
        RECT 53.000 17.900 53.280 18.195 ;
        RECT 48.450 13.445 48.680 17.900 ;
        RECT 50.200 13.800 50.430 17.840 ;
        RECT 49.040 11.700 50.040 11.790 ;
        RECT 48.000 11.560 50.040 11.700 ;
        RECT 48.000 11.500 49.300 11.560 ;
        RECT 49.000 11.300 49.300 11.500 ;
        RECT 49.000 10.800 49.500 11.300 ;
        RECT 50.200 10.600 50.400 13.800 ;
        RECT 50.750 13.445 50.980 17.900 ;
        RECT 52.500 13.800 52.730 17.840 ;
        RECT 51.340 11.560 52.340 11.790 ;
        RECT 51.400 11.300 51.700 11.560 ;
        RECT 51.400 10.800 51.900 11.300 ;
        RECT 52.500 10.600 52.700 13.800 ;
        RECT 53.050 13.700 53.280 17.900 ;
        RECT 54.800 13.800 55.030 17.840 ;
        RECT 53.050 13.445 53.300 13.700 ;
        RECT 53.100 11.300 53.300 13.445 ;
        RECT 53.640 11.560 54.640 11.790 ;
        RECT 53.700 11.300 54.000 11.560 ;
        RECT 53.100 11.100 53.500 11.300 ;
        RECT 50.200 10.100 50.700 10.600 ;
        RECT 52.500 10.100 53.000 10.600 ;
        RECT 53.300 9.900 53.500 11.100 ;
        RECT 53.700 10.800 54.200 11.300 ;
        RECT 54.800 10.600 55.000 13.800 ;
        RECT 54.700 10.100 55.200 10.600 ;
        RECT 55.350 9.900 55.580 16.920 ;
        RECT 53.300 9.700 55.580 9.900 ;
        RECT 54.600 5.500 54.800 9.700 ;
        RECT 55.350 9.620 55.580 9.700 ;
        RECT 57.100 9.975 57.330 16.565 ;
        RECT 57.100 6.700 57.300 9.975 ;
        RECT 58.200 6.700 58.400 21.200 ;
        RECT 69.200 21.000 69.400 23.200 ;
        RECT 65.400 20.950 69.400 21.000 ;
        RECT 60.975 20.800 69.400 20.950 ;
        RECT 60.975 20.720 65.665 20.800 ;
        RECT 69.200 20.400 69.400 20.800 ;
        RECT 66.800 20.380 69.400 20.400 ;
        RECT 59.140 20.200 69.400 20.380 ;
        RECT 59.140 20.150 67.140 20.200 ;
        RECT 67.400 19.890 68.300 19.900 ;
        RECT 67.345 19.400 68.300 19.890 ;
        RECT 67.345 19.350 67.575 19.400 ;
        RECT 59.140 18.860 67.140 19.090 ;
        RECT 59.200 17.985 59.400 18.860 ;
        RECT 69.200 18.600 69.400 20.200 ;
        RECT 65.400 18.555 69.400 18.600 ;
        RECT 60.975 18.400 69.400 18.555 ;
        RECT 60.975 18.325 65.665 18.400 ;
        RECT 59.140 17.755 67.140 17.985 ;
        RECT 67.400 17.495 68.300 17.500 ;
        RECT 67.345 17.000 68.300 17.495 ;
        RECT 67.345 16.955 67.575 17.000 ;
        RECT 59.140 16.600 67.140 16.695 ;
        RECT 68.500 16.600 69.000 16.800 ;
        RECT 59.140 16.465 69.000 16.600 ;
        RECT 66.900 16.400 69.000 16.465 ;
        RECT 68.500 16.300 69.000 16.400 ;
        RECT 69.200 16.100 69.400 18.400 ;
        RECT 62.300 16.050 69.400 16.100 ;
        RECT 62.080 15.900 69.400 16.050 ;
        RECT 62.080 15.820 62.980 15.900 ;
        RECT 59.480 15.500 60.280 15.550 ;
        RECT 56.600 6.690 58.400 6.700 ;
        RECT 55.940 6.500 58.400 6.690 ;
        RECT 58.600 15.320 60.280 15.500 ;
        RECT 62.300 15.480 62.500 15.820 ;
        RECT 63.700 15.550 64.700 15.600 ;
        RECT 58.600 15.300 59.800 15.320 ;
        RECT 58.600 14.900 58.800 15.300 ;
        RECT 62.140 15.250 62.560 15.480 ;
        RECT 63.700 15.400 65.245 15.550 ;
        RECT 59.120 14.900 59.350 14.960 ;
        RECT 58.600 14.700 59.350 14.900 ;
        RECT 55.940 6.460 56.940 6.500 ;
        RECT 56.000 6.200 56.200 6.460 ;
        RECT 56.000 5.700 56.500 6.200 ;
        RECT 58.600 5.500 58.800 14.700 ;
        RECT 59.120 6.960 59.350 14.700 ;
        RECT 60.410 7.300 60.640 14.960 ;
        RECT 62.765 9.500 62.995 13.240 ;
        RECT 62.765 9.200 63.000 9.500 ;
        RECT 60.410 6.960 60.700 7.300 ;
        RECT 62.200 7.190 62.400 7.200 ;
        RECT 62.140 6.960 62.560 7.190 ;
        RECT 59.610 6.570 60.150 6.800 ;
        RECT 59.900 6.300 60.100 6.570 ;
        RECT 59.600 5.800 60.100 6.300 ;
        RECT 60.500 6.300 60.700 6.960 ;
        RECT 60.500 6.000 61.000 6.300 ;
        RECT 62.200 6.000 62.400 6.960 ;
        RECT 60.500 5.800 62.400 6.000 ;
        RECT 54.600 5.300 58.800 5.500 ;
        RECT 59.900 5.600 60.100 5.800 ;
        RECT 62.800 5.600 63.000 9.200 ;
        RECT 59.900 5.400 63.000 5.600 ;
        RECT 63.700 6.700 63.900 15.400 ;
        RECT 64.365 15.320 65.245 15.400 ;
        RECT 67.800 15.000 68.300 15.300 ;
        RECT 64.600 14.980 68.300 15.000 ;
        RECT 64.440 14.800 68.300 14.980 ;
        RECT 68.500 14.800 69.000 15.300 ;
        RECT 64.440 14.750 64.860 14.800 ;
        RECT 68.600 13.100 68.800 14.800 ;
        RECT 65.020 10.700 65.250 12.740 ;
        RECT 65.020 10.500 66.000 10.700 ;
        RECT 65.020 8.700 65.250 10.500 ;
        RECT 65.500 10.200 66.000 10.500 ;
        RECT 67.720 9.400 67.950 13.100 ;
        RECT 67.600 9.100 67.950 9.400 ;
        RECT 68.510 12.800 68.800 13.100 ;
        RECT 68.510 9.100 68.740 12.800 ;
        RECT 69.200 12.265 69.400 15.900 ;
        RECT 69.080 11.900 69.400 12.265 ;
        RECT 69.080 9.575 69.310 11.900 ;
        RECT 63.700 6.690 64.700 6.700 ;
        RECT 63.700 6.500 64.860 6.690 ;
        RECT 58.600 5.200 58.800 5.300 ;
        RECT 63.700 5.200 63.900 6.500 ;
        RECT 64.440 6.460 64.860 6.500 ;
        RECT 58.600 5.000 63.900 5.200 ;
        RECT 67.600 4.800 67.800 9.100 ;
        RECT 68.000 8.665 68.460 8.895 ;
        RECT 68.100 7.900 68.300 8.665 ;
        RECT 68.100 7.200 68.800 7.900 ;
        RECT 68.100 6.200 68.800 6.900 ;
        RECT 71.000 5.000 73.000 42.300 ;
        RECT 73.200 130.800 73.400 168.900 ;
        RECT 86.975 168.500 91.665 168.550 ;
        RECT 97.000 168.500 99.000 210.000 ;
        RECT 74.400 168.000 74.900 168.500 ;
        RECT 86.975 168.320 99.000 168.500 ;
        RECT 91.400 168.300 99.000 168.320 ;
        RECT 82.800 168.000 84.400 168.100 ;
        RECT 95.200 168.000 95.400 168.300 ;
        RECT 74.400 167.640 74.600 168.000 ;
        RECT 75.040 167.900 84.400 168.000 ;
        RECT 92.800 167.980 95.400 168.000 ;
        RECT 75.040 167.770 83.040 167.900 ;
        RECT 74.400 167.500 74.680 167.640 ;
        RECT 74.450 166.840 74.680 167.500 ;
        RECT 83.200 167.500 83.430 167.510 ;
        RECT 83.200 167.000 84.000 167.500 ;
        RECT 83.200 166.970 83.430 167.000 ;
        RECT 75.040 166.600 83.040 166.710 ;
        RECT 74.000 166.480 83.040 166.600 ;
        RECT 74.000 166.400 75.300 166.480 ;
        RECT 74.000 164.200 74.200 166.400 ;
        RECT 74.400 165.500 74.900 166.000 ;
        RECT 84.200 165.600 84.400 167.900 ;
        RECT 85.140 167.800 95.400 167.980 ;
        RECT 85.140 167.750 93.140 167.800 ;
        RECT 93.400 167.490 94.300 167.500 ;
        RECT 93.345 167.000 94.300 167.490 ;
        RECT 93.345 166.950 93.575 167.000 ;
        RECT 85.140 166.460 93.140 166.690 ;
        RECT 82.800 165.570 84.400 165.600 ;
        RECT 74.400 165.210 74.600 165.500 ;
        RECT 75.040 165.400 84.400 165.570 ;
        RECT 85.200 165.550 85.400 166.460 ;
        RECT 86.975 166.100 91.665 166.120 ;
        RECT 95.200 166.100 95.400 167.800 ;
        RECT 86.975 165.900 95.400 166.100 ;
        RECT 86.975 165.890 91.665 165.900 ;
        RECT 75.040 165.340 83.040 165.400 ;
        RECT 74.400 165.000 74.680 165.210 ;
        RECT 83.300 165.080 84.000 165.100 ;
        RECT 74.450 164.410 74.680 165.000 ;
        RECT 83.200 164.600 84.000 165.080 ;
        RECT 83.200 164.540 83.430 164.600 ;
        RECT 75.040 164.200 83.040 164.280 ;
        RECT 74.000 164.050 83.040 164.200 ;
        RECT 74.000 164.000 75.300 164.050 ;
        RECT 74.000 161.800 74.200 164.000 ;
        RECT 74.400 163.100 74.900 163.600 ;
        RECT 84.200 163.200 84.400 165.400 ;
        RECT 85.140 165.320 93.140 165.550 ;
        RECT 93.345 165.000 93.575 165.060 ;
        RECT 93.345 164.520 94.300 165.000 ;
        RECT 93.400 164.500 94.300 164.520 ;
        RECT 85.140 164.030 93.140 164.260 ;
        RECT 82.800 163.140 84.400 163.200 ;
        RECT 74.400 162.780 74.600 163.100 ;
        RECT 75.040 163.000 84.400 163.140 ;
        RECT 75.040 162.910 83.040 163.000 ;
        RECT 74.400 162.600 74.680 162.780 ;
        RECT 83.300 162.650 84.000 162.700 ;
        RECT 74.450 161.980 74.680 162.600 ;
        RECT 83.200 162.200 84.000 162.650 ;
        RECT 83.200 162.110 83.430 162.200 ;
        RECT 75.040 161.800 83.040 161.850 ;
        RECT 74.000 161.620 83.040 161.800 ;
        RECT 74.000 161.600 75.300 161.620 ;
        RECT 74.000 159.300 74.200 161.600 ;
        RECT 74.400 160.700 74.900 161.200 ;
        RECT 84.200 161.100 84.400 163.000 ;
        RECT 85.200 162.580 85.400 164.030 ;
        RECT 86.960 162.920 91.630 163.150 ;
        RECT 91.400 162.900 91.600 162.920 ;
        RECT 92.900 162.580 95.000 162.600 ;
        RECT 85.140 162.400 95.000 162.580 ;
        RECT 85.140 162.350 93.140 162.400 ;
        RECT 93.400 162.090 93.600 162.400 ;
        RECT 94.500 162.100 95.000 162.400 ;
        RECT 93.300 161.900 93.600 162.090 ;
        RECT 93.300 161.550 93.530 161.900 ;
        RECT 85.140 161.200 93.140 161.290 ;
        RECT 84.200 160.800 84.700 161.100 ;
        RECT 82.800 160.710 84.700 160.800 ;
        RECT 74.400 160.350 74.600 160.700 ;
        RECT 75.040 160.600 84.700 160.710 ;
        RECT 84.900 161.060 93.140 161.200 ;
        RECT 84.900 161.000 85.400 161.060 ;
        RECT 75.040 160.480 83.040 160.600 ;
        RECT 84.900 160.400 85.100 161.000 ;
        RECT 74.400 160.100 74.680 160.350 ;
        RECT 74.450 159.550 74.680 160.100 ;
        RECT 83.200 160.200 83.430 160.220 ;
        RECT 84.400 160.200 85.100 160.400 ;
        RECT 95.200 160.200 95.400 165.900 ;
        RECT 83.200 159.700 84.000 160.200 ;
        RECT 83.200 159.680 83.430 159.700 ;
        RECT 75.040 159.300 83.040 159.420 ;
        RECT 74.000 159.190 83.040 159.300 ;
        RECT 74.000 159.100 75.300 159.190 ;
        RECT 74.000 154.500 74.200 159.100 ;
        RECT 74.400 158.300 74.900 158.800 ;
        RECT 84.400 158.300 84.600 160.200 ;
        RECT 91.400 160.150 95.400 160.200 ;
        RECT 86.975 160.000 95.400 160.150 ;
        RECT 86.975 159.920 91.665 160.000 ;
        RECT 95.200 159.600 95.400 160.000 ;
        RECT 92.800 159.580 95.400 159.600 ;
        RECT 85.140 159.400 95.400 159.580 ;
        RECT 85.140 159.350 93.140 159.400 ;
        RECT 93.400 159.090 94.300 159.100 ;
        RECT 93.345 158.600 94.300 159.090 ;
        RECT 93.345 158.550 93.575 158.600 ;
        RECT 74.400 157.920 74.600 158.300 ;
        RECT 82.800 158.280 84.600 158.300 ;
        RECT 75.040 158.100 84.600 158.280 ;
        RECT 75.040 158.050 83.040 158.100 ;
        RECT 74.400 157.120 74.680 157.920 ;
        RECT 83.800 157.800 84.000 158.100 ;
        RECT 85.140 158.060 93.140 158.290 ;
        RECT 83.300 157.790 84.000 157.800 ;
        RECT 83.200 157.300 84.000 157.790 ;
        RECT 83.200 157.250 83.430 157.300 ;
        RECT 85.200 157.150 85.400 158.060 ;
        RECT 86.980 157.700 91.670 157.720 ;
        RECT 95.200 157.700 95.400 159.400 ;
        RECT 86.980 157.500 95.400 157.700 ;
        RECT 86.980 157.490 91.670 157.500 ;
        RECT 74.400 156.900 74.600 157.120 ;
        RECT 75.040 156.900 83.040 156.990 ;
        RECT 85.145 156.920 93.145 157.150 ;
        RECT 74.400 156.760 83.040 156.900 ;
        RECT 74.400 156.700 75.300 156.760 ;
        RECT 93.400 156.660 94.300 156.700 ;
        RECT 74.400 155.800 74.900 156.300 ;
        RECT 93.350 156.200 94.300 156.660 ;
        RECT 84.200 155.900 84.700 156.200 ;
        RECT 93.350 156.120 93.600 156.200 ;
        RECT 82.800 155.850 84.700 155.900 ;
        RECT 74.400 155.490 74.600 155.800 ;
        RECT 75.040 155.700 84.700 155.850 ;
        RECT 75.040 155.620 83.040 155.700 ;
        RECT 74.400 155.300 74.680 155.490 ;
        RECT 74.450 154.690 74.680 155.300 ;
        RECT 83.200 155.300 83.430 155.360 ;
        RECT 83.200 154.820 84.000 155.300 ;
        RECT 83.300 154.800 84.000 154.820 ;
        RECT 75.040 154.500 83.040 154.560 ;
        RECT 74.000 154.330 83.040 154.500 ;
        RECT 74.000 154.300 75.300 154.330 ;
        RECT 74.000 152.100 74.200 154.300 ;
        RECT 74.400 153.400 74.900 153.900 ;
        RECT 84.200 153.500 84.400 155.700 ;
        RECT 85.145 155.630 93.145 155.860 ;
        RECT 85.200 154.170 85.400 155.630 ;
        RECT 86.975 154.510 91.645 154.740 ;
        RECT 93.400 154.200 93.600 156.120 ;
        RECT 92.900 154.170 93.600 154.200 ;
        RECT 85.155 154.000 93.600 154.170 ;
        RECT 85.155 153.940 93.155 154.000 ;
        RECT 94.500 153.700 95.000 153.900 ;
        RECT 93.400 153.680 95.000 153.700 ;
        RECT 82.800 153.420 84.400 153.500 ;
        RECT 74.400 153.060 74.600 153.400 ;
        RECT 75.040 153.300 84.400 153.420 ;
        RECT 75.040 153.190 83.040 153.300 ;
        RECT 74.400 152.900 74.680 153.060 ;
        RECT 74.450 152.260 74.680 152.900 ;
        RECT 83.200 152.900 83.430 152.930 ;
        RECT 83.200 152.400 84.000 152.900 ;
        RECT 84.200 152.800 84.400 153.300 ;
        RECT 93.315 153.400 95.000 153.680 ;
        RECT 93.315 153.140 93.545 153.400 ;
        RECT 85.155 152.800 93.155 152.880 ;
        RECT 84.200 152.650 93.155 152.800 ;
        RECT 84.200 152.600 85.400 152.650 ;
        RECT 83.200 152.390 83.430 152.400 ;
        RECT 75.040 152.100 83.040 152.130 ;
        RECT 74.000 151.900 83.040 152.100 ;
        RECT 74.000 149.600 74.200 151.900 ;
        RECT 74.400 150.900 74.900 151.400 ;
        RECT 84.200 151.000 84.400 152.600 ;
        RECT 95.200 151.800 95.400 157.500 ;
        RECT 91.400 151.750 95.400 151.800 ;
        RECT 86.975 151.600 95.400 151.750 ;
        RECT 86.975 151.520 91.665 151.600 ;
        RECT 95.200 151.200 95.400 151.600 ;
        RECT 92.800 151.180 95.400 151.200 ;
        RECT 82.800 150.990 84.400 151.000 ;
        RECT 74.400 150.630 74.600 150.900 ;
        RECT 75.040 150.800 84.400 150.990 ;
        RECT 85.140 151.000 95.400 151.180 ;
        RECT 85.140 150.950 93.140 151.000 ;
        RECT 75.040 150.760 83.040 150.800 ;
        RECT 74.400 150.400 74.680 150.630 ;
        RECT 74.450 149.830 74.680 150.400 ;
        RECT 83.200 150.000 84.000 150.500 ;
        RECT 83.200 149.960 83.430 150.000 ;
        RECT 75.040 149.600 83.040 149.700 ;
        RECT 74.000 149.470 83.040 149.600 ;
        RECT 74.000 149.400 75.300 149.470 ;
        RECT 74.000 147.200 74.200 149.400 ;
        RECT 74.400 148.500 74.900 149.000 ;
        RECT 84.200 148.600 84.400 150.800 ;
        RECT 93.400 150.690 94.300 150.700 ;
        RECT 93.345 150.200 94.300 150.690 ;
        RECT 93.345 150.150 93.575 150.200 ;
        RECT 85.140 149.660 93.140 149.890 ;
        RECT 85.300 148.780 85.500 149.660 ;
        RECT 95.200 149.400 95.400 151.000 ;
        RECT 91.400 149.350 95.400 149.400 ;
        RECT 86.975 149.200 95.400 149.350 ;
        RECT 86.975 149.120 91.665 149.200 ;
        RECT 82.800 148.560 84.400 148.600 ;
        RECT 74.400 148.200 74.600 148.500 ;
        RECT 75.040 148.400 84.400 148.560 ;
        RECT 85.140 148.550 93.140 148.780 ;
        RECT 75.040 148.330 83.040 148.400 ;
        RECT 93.400 148.290 94.300 148.300 ;
        RECT 74.400 147.900 74.680 148.200 ;
        RECT 83.300 148.070 84.000 148.100 ;
        RECT 74.450 147.400 74.680 147.900 ;
        RECT 83.200 147.600 84.000 148.070 ;
        RECT 93.345 147.800 94.300 148.290 ;
        RECT 93.345 147.750 93.575 147.800 ;
        RECT 83.200 147.530 83.430 147.600 ;
        RECT 85.140 147.400 93.140 147.490 ;
        RECT 75.040 147.200 83.040 147.270 ;
        RECT 74.000 147.040 83.040 147.200 ;
        RECT 84.200 147.260 93.140 147.400 ;
        RECT 84.200 147.200 85.400 147.260 ;
        RECT 74.000 147.000 75.300 147.040 ;
        RECT 74.000 137.700 74.200 147.000 ;
        RECT 74.400 146.500 79.200 146.700 ;
        RECT 74.400 146.100 74.900 146.500 ;
        RECT 76.700 146.100 76.900 146.500 ;
        RECT 74.400 146.080 75.400 146.100 ;
        RECT 76.700 146.080 77.700 146.100 ;
        RECT 74.400 145.900 76.040 146.080 ;
        RECT 74.400 144.195 74.600 145.900 ;
        RECT 75.040 145.850 76.040 145.900 ;
        RECT 76.700 145.900 78.340 146.080 ;
        RECT 76.700 144.195 76.900 145.900 ;
        RECT 77.340 145.850 78.340 145.900 ;
        RECT 79.000 144.195 79.200 146.500 ;
        RECT 80.300 146.080 82.200 146.100 ;
        RECT 79.640 145.900 82.940 146.080 ;
        RECT 79.640 145.850 80.640 145.900 ;
        RECT 81.940 145.850 82.940 145.900 ;
        RECT 74.400 143.900 74.680 144.195 ;
        RECT 76.700 143.900 76.980 144.195 ;
        RECT 79.000 143.900 79.280 144.195 ;
        RECT 74.450 139.445 74.680 143.900 ;
        RECT 76.200 139.800 76.430 143.840 ;
        RECT 75.040 137.700 76.040 137.790 ;
        RECT 74.000 137.560 76.040 137.700 ;
        RECT 74.000 137.500 75.300 137.560 ;
        RECT 75.000 137.300 75.300 137.500 ;
        RECT 75.000 136.800 75.500 137.300 ;
        RECT 76.200 136.600 76.400 139.800 ;
        RECT 76.750 139.445 76.980 143.900 ;
        RECT 78.500 139.800 78.730 143.840 ;
        RECT 77.340 137.560 78.340 137.790 ;
        RECT 77.400 137.300 77.700 137.560 ;
        RECT 77.400 136.800 77.900 137.300 ;
        RECT 78.500 136.600 78.700 139.800 ;
        RECT 79.050 139.700 79.280 143.900 ;
        RECT 80.800 139.800 81.030 143.840 ;
        RECT 79.050 139.445 79.300 139.700 ;
        RECT 79.100 137.300 79.300 139.445 ;
        RECT 79.640 137.560 80.640 137.790 ;
        RECT 79.700 137.300 80.000 137.560 ;
        RECT 79.100 137.100 79.500 137.300 ;
        RECT 76.200 136.100 76.700 136.600 ;
        RECT 78.500 136.100 79.000 136.600 ;
        RECT 79.300 135.900 79.500 137.100 ;
        RECT 79.700 136.800 80.200 137.300 ;
        RECT 80.800 136.600 81.000 139.800 ;
        RECT 80.700 136.100 81.200 136.600 ;
        RECT 81.350 135.900 81.580 142.920 ;
        RECT 79.300 135.700 81.580 135.900 ;
        RECT 80.600 131.500 80.800 135.700 ;
        RECT 81.350 135.620 81.580 135.700 ;
        RECT 83.100 135.975 83.330 142.565 ;
        RECT 83.100 132.700 83.300 135.975 ;
        RECT 84.200 132.700 84.400 147.200 ;
        RECT 95.200 147.000 95.400 149.200 ;
        RECT 91.400 146.950 95.400 147.000 ;
        RECT 86.975 146.800 95.400 146.950 ;
        RECT 86.975 146.720 91.665 146.800 ;
        RECT 95.200 146.400 95.400 146.800 ;
        RECT 92.800 146.380 95.400 146.400 ;
        RECT 85.140 146.200 95.400 146.380 ;
        RECT 85.140 146.150 93.140 146.200 ;
        RECT 93.400 145.890 94.300 145.900 ;
        RECT 93.345 145.400 94.300 145.890 ;
        RECT 93.345 145.350 93.575 145.400 ;
        RECT 85.140 144.860 93.140 145.090 ;
        RECT 85.200 143.985 85.400 144.860 ;
        RECT 95.200 144.600 95.400 146.200 ;
        RECT 91.400 144.555 95.400 144.600 ;
        RECT 86.975 144.400 95.400 144.555 ;
        RECT 86.975 144.325 91.665 144.400 ;
        RECT 85.140 143.755 93.140 143.985 ;
        RECT 93.400 143.495 94.300 143.500 ;
        RECT 93.345 143.000 94.300 143.495 ;
        RECT 93.345 142.955 93.575 143.000 ;
        RECT 85.140 142.600 93.140 142.695 ;
        RECT 94.500 142.600 95.000 142.800 ;
        RECT 85.140 142.465 95.000 142.600 ;
        RECT 92.900 142.400 95.000 142.465 ;
        RECT 94.500 142.300 95.000 142.400 ;
        RECT 95.200 142.100 95.400 144.400 ;
        RECT 88.300 142.050 95.400 142.100 ;
        RECT 88.080 141.900 95.400 142.050 ;
        RECT 88.080 141.820 88.980 141.900 ;
        RECT 85.480 141.500 86.280 141.550 ;
        RECT 82.600 132.690 84.400 132.700 ;
        RECT 81.940 132.500 84.400 132.690 ;
        RECT 84.600 141.320 86.280 141.500 ;
        RECT 88.300 141.480 88.500 141.820 ;
        RECT 89.700 141.550 90.700 141.600 ;
        RECT 84.600 141.300 85.800 141.320 ;
        RECT 84.600 140.900 84.800 141.300 ;
        RECT 88.140 141.250 88.560 141.480 ;
        RECT 89.700 141.400 91.245 141.550 ;
        RECT 85.120 140.900 85.350 140.960 ;
        RECT 84.600 140.700 85.350 140.900 ;
        RECT 81.940 132.460 82.940 132.500 ;
        RECT 82.000 132.200 82.200 132.460 ;
        RECT 82.000 131.700 82.500 132.200 ;
        RECT 84.600 131.500 84.800 140.700 ;
        RECT 85.120 132.960 85.350 140.700 ;
        RECT 86.410 133.300 86.640 140.960 ;
        RECT 88.765 135.500 88.995 139.240 ;
        RECT 88.765 135.200 89.000 135.500 ;
        RECT 86.410 132.960 86.700 133.300 ;
        RECT 88.200 133.190 88.400 133.200 ;
        RECT 88.140 132.960 88.560 133.190 ;
        RECT 85.610 132.570 86.150 132.800 ;
        RECT 85.900 132.300 86.100 132.570 ;
        RECT 85.600 131.800 86.100 132.300 ;
        RECT 86.500 132.300 86.700 132.960 ;
        RECT 86.500 132.000 87.000 132.300 ;
        RECT 88.200 132.000 88.400 132.960 ;
        RECT 86.500 131.800 88.400 132.000 ;
        RECT 80.600 131.300 84.800 131.500 ;
        RECT 85.900 131.600 86.100 131.800 ;
        RECT 88.800 131.600 89.000 135.200 ;
        RECT 85.900 131.400 89.000 131.600 ;
        RECT 89.700 132.700 89.900 141.400 ;
        RECT 90.365 141.320 91.245 141.400 ;
        RECT 93.800 141.000 94.300 141.300 ;
        RECT 90.600 140.980 94.300 141.000 ;
        RECT 90.440 140.800 94.300 140.980 ;
        RECT 94.500 140.800 95.000 141.300 ;
        RECT 90.440 140.750 90.860 140.800 ;
        RECT 94.600 139.100 94.800 140.800 ;
        RECT 91.020 136.700 91.250 138.740 ;
        RECT 91.020 136.500 92.000 136.700 ;
        RECT 91.020 134.700 91.250 136.500 ;
        RECT 91.500 136.200 92.000 136.500 ;
        RECT 93.720 135.400 93.950 139.100 ;
        RECT 93.600 135.100 93.950 135.400 ;
        RECT 94.510 138.800 94.800 139.100 ;
        RECT 94.510 135.100 94.740 138.800 ;
        RECT 95.200 138.265 95.400 141.900 ;
        RECT 95.080 138.000 95.400 138.265 ;
        RECT 95.080 135.575 95.310 138.000 ;
        RECT 89.700 132.690 90.700 132.700 ;
        RECT 89.700 132.500 90.860 132.690 ;
        RECT 84.600 131.200 84.800 131.300 ;
        RECT 89.700 131.200 89.900 132.500 ;
        RECT 90.440 132.460 90.860 132.500 ;
        RECT 84.600 131.000 89.900 131.200 ;
        RECT 93.600 130.800 93.800 135.100 ;
        RECT 94.000 134.665 94.460 134.895 ;
        RECT 94.100 133.900 94.300 134.665 ;
        RECT 94.100 133.200 94.800 133.900 ;
        RECT 94.100 132.200 94.800 132.900 ;
        RECT 73.200 130.600 93.800 130.800 ;
        RECT 73.200 88.800 73.400 130.600 ;
        RECT 86.975 126.500 91.665 126.550 ;
        RECT 97.000 126.500 99.000 168.300 ;
        RECT 74.400 126.000 74.900 126.500 ;
        RECT 86.975 126.320 99.000 126.500 ;
        RECT 91.400 126.300 99.000 126.320 ;
        RECT 82.800 126.000 84.400 126.100 ;
        RECT 95.200 126.000 95.400 126.300 ;
        RECT 74.400 125.640 74.600 126.000 ;
        RECT 75.040 125.900 84.400 126.000 ;
        RECT 92.800 125.980 95.400 126.000 ;
        RECT 75.040 125.770 83.040 125.900 ;
        RECT 74.400 125.500 74.680 125.640 ;
        RECT 74.450 124.840 74.680 125.500 ;
        RECT 83.200 125.500 83.430 125.510 ;
        RECT 83.200 125.000 84.000 125.500 ;
        RECT 83.200 124.970 83.430 125.000 ;
        RECT 75.040 124.600 83.040 124.710 ;
        RECT 74.000 124.480 83.040 124.600 ;
        RECT 74.000 124.400 75.300 124.480 ;
        RECT 74.000 122.200 74.200 124.400 ;
        RECT 74.400 123.500 74.900 124.000 ;
        RECT 84.200 123.600 84.400 125.900 ;
        RECT 85.140 125.800 95.400 125.980 ;
        RECT 85.140 125.750 93.140 125.800 ;
        RECT 93.400 125.490 94.300 125.500 ;
        RECT 93.345 125.000 94.300 125.490 ;
        RECT 93.345 124.950 93.575 125.000 ;
        RECT 85.140 124.460 93.140 124.690 ;
        RECT 82.800 123.570 84.400 123.600 ;
        RECT 74.400 123.210 74.600 123.500 ;
        RECT 75.040 123.400 84.400 123.570 ;
        RECT 85.200 123.550 85.400 124.460 ;
        RECT 86.975 124.100 91.665 124.120 ;
        RECT 95.200 124.100 95.400 125.800 ;
        RECT 86.975 123.900 95.400 124.100 ;
        RECT 86.975 123.890 91.665 123.900 ;
        RECT 75.040 123.340 83.040 123.400 ;
        RECT 74.400 123.000 74.680 123.210 ;
        RECT 83.300 123.080 84.000 123.100 ;
        RECT 74.450 122.410 74.680 123.000 ;
        RECT 83.200 122.600 84.000 123.080 ;
        RECT 83.200 122.540 83.430 122.600 ;
        RECT 75.040 122.200 83.040 122.280 ;
        RECT 74.000 122.050 83.040 122.200 ;
        RECT 74.000 122.000 75.300 122.050 ;
        RECT 74.000 119.800 74.200 122.000 ;
        RECT 74.400 121.100 74.900 121.600 ;
        RECT 84.200 121.200 84.400 123.400 ;
        RECT 85.140 123.320 93.140 123.550 ;
        RECT 93.345 123.000 93.575 123.060 ;
        RECT 93.345 122.520 94.300 123.000 ;
        RECT 93.400 122.500 94.300 122.520 ;
        RECT 85.140 122.030 93.140 122.260 ;
        RECT 82.800 121.140 84.400 121.200 ;
        RECT 74.400 120.780 74.600 121.100 ;
        RECT 75.040 121.000 84.400 121.140 ;
        RECT 75.040 120.910 83.040 121.000 ;
        RECT 74.400 120.600 74.680 120.780 ;
        RECT 83.300 120.650 84.000 120.700 ;
        RECT 74.450 119.980 74.680 120.600 ;
        RECT 83.200 120.200 84.000 120.650 ;
        RECT 83.200 120.110 83.430 120.200 ;
        RECT 75.040 119.800 83.040 119.850 ;
        RECT 74.000 119.620 83.040 119.800 ;
        RECT 74.000 119.600 75.300 119.620 ;
        RECT 74.000 117.300 74.200 119.600 ;
        RECT 74.400 118.700 74.900 119.200 ;
        RECT 84.200 119.100 84.400 121.000 ;
        RECT 85.200 120.580 85.400 122.030 ;
        RECT 86.960 120.920 91.630 121.150 ;
        RECT 91.400 120.900 91.600 120.920 ;
        RECT 92.900 120.580 95.000 120.600 ;
        RECT 85.140 120.400 95.000 120.580 ;
        RECT 85.140 120.350 93.140 120.400 ;
        RECT 93.400 120.090 93.600 120.400 ;
        RECT 94.500 120.100 95.000 120.400 ;
        RECT 93.300 119.900 93.600 120.090 ;
        RECT 93.300 119.550 93.530 119.900 ;
        RECT 85.140 119.200 93.140 119.290 ;
        RECT 84.200 118.800 84.700 119.100 ;
        RECT 82.800 118.710 84.700 118.800 ;
        RECT 74.400 118.350 74.600 118.700 ;
        RECT 75.040 118.600 84.700 118.710 ;
        RECT 84.900 119.060 93.140 119.200 ;
        RECT 84.900 119.000 85.400 119.060 ;
        RECT 75.040 118.480 83.040 118.600 ;
        RECT 84.900 118.400 85.100 119.000 ;
        RECT 74.400 118.100 74.680 118.350 ;
        RECT 74.450 117.550 74.680 118.100 ;
        RECT 83.200 118.200 83.430 118.220 ;
        RECT 84.400 118.200 85.100 118.400 ;
        RECT 95.200 118.200 95.400 123.900 ;
        RECT 83.200 117.700 84.000 118.200 ;
        RECT 83.200 117.680 83.430 117.700 ;
        RECT 75.040 117.300 83.040 117.420 ;
        RECT 74.000 117.190 83.040 117.300 ;
        RECT 74.000 117.100 75.300 117.190 ;
        RECT 74.000 112.500 74.200 117.100 ;
        RECT 74.400 116.300 74.900 116.800 ;
        RECT 84.400 116.300 84.600 118.200 ;
        RECT 91.400 118.150 95.400 118.200 ;
        RECT 86.975 118.000 95.400 118.150 ;
        RECT 86.975 117.920 91.665 118.000 ;
        RECT 95.200 117.600 95.400 118.000 ;
        RECT 92.800 117.580 95.400 117.600 ;
        RECT 85.140 117.400 95.400 117.580 ;
        RECT 85.140 117.350 93.140 117.400 ;
        RECT 93.400 117.090 94.300 117.100 ;
        RECT 93.345 116.600 94.300 117.090 ;
        RECT 93.345 116.550 93.575 116.600 ;
        RECT 74.400 115.920 74.600 116.300 ;
        RECT 82.800 116.280 84.600 116.300 ;
        RECT 75.040 116.100 84.600 116.280 ;
        RECT 75.040 116.050 83.040 116.100 ;
        RECT 74.400 115.120 74.680 115.920 ;
        RECT 83.800 115.800 84.000 116.100 ;
        RECT 85.140 116.060 93.140 116.290 ;
        RECT 83.300 115.790 84.000 115.800 ;
        RECT 83.200 115.300 84.000 115.790 ;
        RECT 83.200 115.250 83.430 115.300 ;
        RECT 85.200 115.150 85.400 116.060 ;
        RECT 86.980 115.700 91.670 115.720 ;
        RECT 95.200 115.700 95.400 117.400 ;
        RECT 86.980 115.500 95.400 115.700 ;
        RECT 86.980 115.490 91.670 115.500 ;
        RECT 74.400 114.900 74.600 115.120 ;
        RECT 75.040 114.900 83.040 114.990 ;
        RECT 85.145 114.920 93.145 115.150 ;
        RECT 74.400 114.760 83.040 114.900 ;
        RECT 74.400 114.700 75.300 114.760 ;
        RECT 93.400 114.660 94.300 114.700 ;
        RECT 74.400 113.800 74.900 114.300 ;
        RECT 93.350 114.200 94.300 114.660 ;
        RECT 84.200 113.900 84.700 114.200 ;
        RECT 93.350 114.120 93.600 114.200 ;
        RECT 82.800 113.850 84.700 113.900 ;
        RECT 74.400 113.490 74.600 113.800 ;
        RECT 75.040 113.700 84.700 113.850 ;
        RECT 75.040 113.620 83.040 113.700 ;
        RECT 74.400 113.300 74.680 113.490 ;
        RECT 74.450 112.690 74.680 113.300 ;
        RECT 83.200 113.300 83.430 113.360 ;
        RECT 83.200 112.820 84.000 113.300 ;
        RECT 83.300 112.800 84.000 112.820 ;
        RECT 75.040 112.500 83.040 112.560 ;
        RECT 74.000 112.330 83.040 112.500 ;
        RECT 74.000 112.300 75.300 112.330 ;
        RECT 74.000 110.100 74.200 112.300 ;
        RECT 74.400 111.400 74.900 111.900 ;
        RECT 84.200 111.500 84.400 113.700 ;
        RECT 85.145 113.630 93.145 113.860 ;
        RECT 85.200 112.170 85.400 113.630 ;
        RECT 86.975 112.510 91.645 112.740 ;
        RECT 93.400 112.200 93.600 114.120 ;
        RECT 92.900 112.170 93.600 112.200 ;
        RECT 85.155 112.000 93.600 112.170 ;
        RECT 85.155 111.940 93.155 112.000 ;
        RECT 94.500 111.700 95.000 111.900 ;
        RECT 93.400 111.680 95.000 111.700 ;
        RECT 82.800 111.420 84.400 111.500 ;
        RECT 74.400 111.060 74.600 111.400 ;
        RECT 75.040 111.300 84.400 111.420 ;
        RECT 75.040 111.190 83.040 111.300 ;
        RECT 74.400 110.900 74.680 111.060 ;
        RECT 74.450 110.260 74.680 110.900 ;
        RECT 83.200 110.900 83.430 110.930 ;
        RECT 83.200 110.400 84.000 110.900 ;
        RECT 84.200 110.800 84.400 111.300 ;
        RECT 93.315 111.400 95.000 111.680 ;
        RECT 93.315 111.140 93.545 111.400 ;
        RECT 85.155 110.800 93.155 110.880 ;
        RECT 84.200 110.650 93.155 110.800 ;
        RECT 84.200 110.600 85.400 110.650 ;
        RECT 83.200 110.390 83.430 110.400 ;
        RECT 75.040 110.100 83.040 110.130 ;
        RECT 74.000 109.900 83.040 110.100 ;
        RECT 74.000 107.600 74.200 109.900 ;
        RECT 74.400 108.900 74.900 109.400 ;
        RECT 84.200 109.000 84.400 110.600 ;
        RECT 95.200 109.800 95.400 115.500 ;
        RECT 91.400 109.750 95.400 109.800 ;
        RECT 86.975 109.600 95.400 109.750 ;
        RECT 86.975 109.520 91.665 109.600 ;
        RECT 95.200 109.200 95.400 109.600 ;
        RECT 92.800 109.180 95.400 109.200 ;
        RECT 82.800 108.990 84.400 109.000 ;
        RECT 74.400 108.630 74.600 108.900 ;
        RECT 75.040 108.800 84.400 108.990 ;
        RECT 85.140 109.000 95.400 109.180 ;
        RECT 85.140 108.950 93.140 109.000 ;
        RECT 75.040 108.760 83.040 108.800 ;
        RECT 74.400 108.400 74.680 108.630 ;
        RECT 74.450 107.830 74.680 108.400 ;
        RECT 83.200 108.000 84.000 108.500 ;
        RECT 83.200 107.960 83.430 108.000 ;
        RECT 75.040 107.600 83.040 107.700 ;
        RECT 74.000 107.470 83.040 107.600 ;
        RECT 74.000 107.400 75.300 107.470 ;
        RECT 74.000 105.200 74.200 107.400 ;
        RECT 74.400 106.500 74.900 107.000 ;
        RECT 84.200 106.600 84.400 108.800 ;
        RECT 93.400 108.690 94.300 108.700 ;
        RECT 93.345 108.200 94.300 108.690 ;
        RECT 93.345 108.150 93.575 108.200 ;
        RECT 85.140 107.660 93.140 107.890 ;
        RECT 85.300 106.780 85.500 107.660 ;
        RECT 95.200 107.400 95.400 109.000 ;
        RECT 91.400 107.350 95.400 107.400 ;
        RECT 86.975 107.200 95.400 107.350 ;
        RECT 86.975 107.120 91.665 107.200 ;
        RECT 82.800 106.560 84.400 106.600 ;
        RECT 74.400 106.200 74.600 106.500 ;
        RECT 75.040 106.400 84.400 106.560 ;
        RECT 85.140 106.550 93.140 106.780 ;
        RECT 75.040 106.330 83.040 106.400 ;
        RECT 93.400 106.290 94.300 106.300 ;
        RECT 74.400 105.900 74.680 106.200 ;
        RECT 83.300 106.070 84.000 106.100 ;
        RECT 74.450 105.400 74.680 105.900 ;
        RECT 83.200 105.600 84.000 106.070 ;
        RECT 93.345 105.800 94.300 106.290 ;
        RECT 93.345 105.750 93.575 105.800 ;
        RECT 83.200 105.530 83.430 105.600 ;
        RECT 85.140 105.400 93.140 105.490 ;
        RECT 75.040 105.200 83.040 105.270 ;
        RECT 74.000 105.040 83.040 105.200 ;
        RECT 84.200 105.260 93.140 105.400 ;
        RECT 84.200 105.200 85.400 105.260 ;
        RECT 74.000 105.000 75.300 105.040 ;
        RECT 74.000 95.700 74.200 105.000 ;
        RECT 74.400 104.500 79.200 104.700 ;
        RECT 74.400 104.100 74.900 104.500 ;
        RECT 76.700 104.100 76.900 104.500 ;
        RECT 74.400 104.080 75.400 104.100 ;
        RECT 76.700 104.080 77.700 104.100 ;
        RECT 74.400 103.900 76.040 104.080 ;
        RECT 74.400 102.195 74.600 103.900 ;
        RECT 75.040 103.850 76.040 103.900 ;
        RECT 76.700 103.900 78.340 104.080 ;
        RECT 76.700 102.195 76.900 103.900 ;
        RECT 77.340 103.850 78.340 103.900 ;
        RECT 79.000 102.195 79.200 104.500 ;
        RECT 80.300 104.080 82.200 104.100 ;
        RECT 79.640 103.900 82.940 104.080 ;
        RECT 79.640 103.850 80.640 103.900 ;
        RECT 81.940 103.850 82.940 103.900 ;
        RECT 74.400 101.900 74.680 102.195 ;
        RECT 76.700 101.900 76.980 102.195 ;
        RECT 79.000 101.900 79.280 102.195 ;
        RECT 74.450 97.445 74.680 101.900 ;
        RECT 76.200 97.800 76.430 101.840 ;
        RECT 75.040 95.700 76.040 95.790 ;
        RECT 74.000 95.560 76.040 95.700 ;
        RECT 74.000 95.500 75.300 95.560 ;
        RECT 75.000 95.300 75.300 95.500 ;
        RECT 75.000 94.800 75.500 95.300 ;
        RECT 76.200 94.600 76.400 97.800 ;
        RECT 76.750 97.445 76.980 101.900 ;
        RECT 78.500 97.800 78.730 101.840 ;
        RECT 77.340 95.560 78.340 95.790 ;
        RECT 77.400 95.300 77.700 95.560 ;
        RECT 77.400 94.800 77.900 95.300 ;
        RECT 78.500 94.600 78.700 97.800 ;
        RECT 79.050 97.700 79.280 101.900 ;
        RECT 80.800 97.800 81.030 101.840 ;
        RECT 79.050 97.445 79.300 97.700 ;
        RECT 79.100 95.300 79.300 97.445 ;
        RECT 79.640 95.560 80.640 95.790 ;
        RECT 79.700 95.300 80.000 95.560 ;
        RECT 79.100 95.100 79.500 95.300 ;
        RECT 76.200 94.100 76.700 94.600 ;
        RECT 78.500 94.100 79.000 94.600 ;
        RECT 79.300 93.900 79.500 95.100 ;
        RECT 79.700 94.800 80.200 95.300 ;
        RECT 80.800 94.600 81.000 97.800 ;
        RECT 80.700 94.100 81.200 94.600 ;
        RECT 81.350 93.900 81.580 100.920 ;
        RECT 79.300 93.700 81.580 93.900 ;
        RECT 80.600 89.500 80.800 93.700 ;
        RECT 81.350 93.620 81.580 93.700 ;
        RECT 83.100 93.975 83.330 100.565 ;
        RECT 83.100 90.700 83.300 93.975 ;
        RECT 84.200 90.700 84.400 105.200 ;
        RECT 95.200 105.000 95.400 107.200 ;
        RECT 91.400 104.950 95.400 105.000 ;
        RECT 86.975 104.800 95.400 104.950 ;
        RECT 86.975 104.720 91.665 104.800 ;
        RECT 95.200 104.400 95.400 104.800 ;
        RECT 92.800 104.380 95.400 104.400 ;
        RECT 85.140 104.200 95.400 104.380 ;
        RECT 85.140 104.150 93.140 104.200 ;
        RECT 93.400 103.890 94.300 103.900 ;
        RECT 93.345 103.400 94.300 103.890 ;
        RECT 93.345 103.350 93.575 103.400 ;
        RECT 85.140 102.860 93.140 103.090 ;
        RECT 85.200 101.985 85.400 102.860 ;
        RECT 95.200 102.600 95.400 104.200 ;
        RECT 91.400 102.555 95.400 102.600 ;
        RECT 86.975 102.400 95.400 102.555 ;
        RECT 86.975 102.325 91.665 102.400 ;
        RECT 85.140 101.755 93.140 101.985 ;
        RECT 93.400 101.495 94.300 101.500 ;
        RECT 93.345 101.000 94.300 101.495 ;
        RECT 93.345 100.955 93.575 101.000 ;
        RECT 85.140 100.600 93.140 100.695 ;
        RECT 94.500 100.600 95.000 100.800 ;
        RECT 85.140 100.465 95.000 100.600 ;
        RECT 92.900 100.400 95.000 100.465 ;
        RECT 94.500 100.300 95.000 100.400 ;
        RECT 95.200 100.100 95.400 102.400 ;
        RECT 88.300 100.050 95.400 100.100 ;
        RECT 88.080 99.900 95.400 100.050 ;
        RECT 88.080 99.820 88.980 99.900 ;
        RECT 85.480 99.500 86.280 99.550 ;
        RECT 82.600 90.690 84.400 90.700 ;
        RECT 81.940 90.500 84.400 90.690 ;
        RECT 84.600 99.320 86.280 99.500 ;
        RECT 88.300 99.480 88.500 99.820 ;
        RECT 89.700 99.550 90.700 99.600 ;
        RECT 84.600 99.300 85.800 99.320 ;
        RECT 84.600 98.900 84.800 99.300 ;
        RECT 88.140 99.250 88.560 99.480 ;
        RECT 89.700 99.400 91.245 99.550 ;
        RECT 85.120 98.900 85.350 98.960 ;
        RECT 84.600 98.700 85.350 98.900 ;
        RECT 81.940 90.460 82.940 90.500 ;
        RECT 82.000 90.200 82.200 90.460 ;
        RECT 82.000 89.700 82.500 90.200 ;
        RECT 84.600 89.500 84.800 98.700 ;
        RECT 85.120 90.960 85.350 98.700 ;
        RECT 86.410 91.300 86.640 98.960 ;
        RECT 88.765 93.500 88.995 97.240 ;
        RECT 88.765 93.200 89.000 93.500 ;
        RECT 86.410 90.960 86.700 91.300 ;
        RECT 88.200 91.190 88.400 91.200 ;
        RECT 88.140 90.960 88.560 91.190 ;
        RECT 85.610 90.570 86.150 90.800 ;
        RECT 85.900 90.300 86.100 90.570 ;
        RECT 85.600 89.800 86.100 90.300 ;
        RECT 86.500 90.300 86.700 90.960 ;
        RECT 86.500 90.000 87.000 90.300 ;
        RECT 88.200 90.000 88.400 90.960 ;
        RECT 86.500 89.800 88.400 90.000 ;
        RECT 80.600 89.300 84.800 89.500 ;
        RECT 85.900 89.600 86.100 89.800 ;
        RECT 88.800 89.600 89.000 93.200 ;
        RECT 85.900 89.400 89.000 89.600 ;
        RECT 89.700 90.700 89.900 99.400 ;
        RECT 90.365 99.320 91.245 99.400 ;
        RECT 93.800 99.000 94.300 99.300 ;
        RECT 90.600 98.980 94.300 99.000 ;
        RECT 90.440 98.800 94.300 98.980 ;
        RECT 94.500 98.800 95.000 99.300 ;
        RECT 90.440 98.750 90.860 98.800 ;
        RECT 94.600 97.100 94.800 98.800 ;
        RECT 91.020 94.700 91.250 96.740 ;
        RECT 91.020 94.500 92.000 94.700 ;
        RECT 91.020 92.700 91.250 94.500 ;
        RECT 91.500 94.200 92.000 94.500 ;
        RECT 93.720 93.400 93.950 97.100 ;
        RECT 93.600 93.100 93.950 93.400 ;
        RECT 94.510 96.800 94.800 97.100 ;
        RECT 94.510 93.100 94.740 96.800 ;
        RECT 95.200 96.265 95.400 99.900 ;
        RECT 95.080 96.000 95.400 96.265 ;
        RECT 95.080 93.575 95.310 96.000 ;
        RECT 89.700 90.690 90.700 90.700 ;
        RECT 89.700 90.500 90.860 90.690 ;
        RECT 84.600 89.200 84.800 89.300 ;
        RECT 89.700 89.200 89.900 90.500 ;
        RECT 90.440 90.460 90.860 90.500 ;
        RECT 84.600 89.000 89.900 89.200 ;
        RECT 93.600 88.800 93.800 93.100 ;
        RECT 94.000 92.665 94.460 92.895 ;
        RECT 94.100 91.900 94.300 92.665 ;
        RECT 94.100 91.200 94.800 91.900 ;
        RECT 94.100 90.200 94.800 90.900 ;
        RECT 73.200 88.600 93.800 88.800 ;
        RECT 73.200 46.800 73.400 88.600 ;
        RECT 86.975 84.500 91.665 84.550 ;
        RECT 97.000 84.500 99.000 126.300 ;
        RECT 74.400 84.000 74.900 84.500 ;
        RECT 86.975 84.320 99.000 84.500 ;
        RECT 91.400 84.300 99.000 84.320 ;
        RECT 82.800 84.000 84.400 84.100 ;
        RECT 95.200 84.000 95.400 84.300 ;
        RECT 74.400 83.640 74.600 84.000 ;
        RECT 75.040 83.900 84.400 84.000 ;
        RECT 92.800 83.980 95.400 84.000 ;
        RECT 75.040 83.770 83.040 83.900 ;
        RECT 74.400 83.500 74.680 83.640 ;
        RECT 74.450 82.840 74.680 83.500 ;
        RECT 83.200 83.500 83.430 83.510 ;
        RECT 83.200 83.000 84.000 83.500 ;
        RECT 83.200 82.970 83.430 83.000 ;
        RECT 75.040 82.600 83.040 82.710 ;
        RECT 74.000 82.480 83.040 82.600 ;
        RECT 74.000 82.400 75.300 82.480 ;
        RECT 74.000 80.200 74.200 82.400 ;
        RECT 74.400 81.500 74.900 82.000 ;
        RECT 84.200 81.600 84.400 83.900 ;
        RECT 85.140 83.800 95.400 83.980 ;
        RECT 85.140 83.750 93.140 83.800 ;
        RECT 93.400 83.490 94.300 83.500 ;
        RECT 93.345 83.000 94.300 83.490 ;
        RECT 93.345 82.950 93.575 83.000 ;
        RECT 85.140 82.460 93.140 82.690 ;
        RECT 82.800 81.570 84.400 81.600 ;
        RECT 74.400 81.210 74.600 81.500 ;
        RECT 75.040 81.400 84.400 81.570 ;
        RECT 85.200 81.550 85.400 82.460 ;
        RECT 86.975 82.100 91.665 82.120 ;
        RECT 95.200 82.100 95.400 83.800 ;
        RECT 86.975 81.900 95.400 82.100 ;
        RECT 86.975 81.890 91.665 81.900 ;
        RECT 75.040 81.340 83.040 81.400 ;
        RECT 74.400 81.000 74.680 81.210 ;
        RECT 83.300 81.080 84.000 81.100 ;
        RECT 74.450 80.410 74.680 81.000 ;
        RECT 83.200 80.600 84.000 81.080 ;
        RECT 83.200 80.540 83.430 80.600 ;
        RECT 75.040 80.200 83.040 80.280 ;
        RECT 74.000 80.050 83.040 80.200 ;
        RECT 74.000 80.000 75.300 80.050 ;
        RECT 74.000 77.800 74.200 80.000 ;
        RECT 74.400 79.100 74.900 79.600 ;
        RECT 84.200 79.200 84.400 81.400 ;
        RECT 85.140 81.320 93.140 81.550 ;
        RECT 93.345 81.000 93.575 81.060 ;
        RECT 93.345 80.520 94.300 81.000 ;
        RECT 93.400 80.500 94.300 80.520 ;
        RECT 85.140 80.030 93.140 80.260 ;
        RECT 82.800 79.140 84.400 79.200 ;
        RECT 74.400 78.780 74.600 79.100 ;
        RECT 75.040 79.000 84.400 79.140 ;
        RECT 75.040 78.910 83.040 79.000 ;
        RECT 74.400 78.600 74.680 78.780 ;
        RECT 83.300 78.650 84.000 78.700 ;
        RECT 74.450 77.980 74.680 78.600 ;
        RECT 83.200 78.200 84.000 78.650 ;
        RECT 83.200 78.110 83.430 78.200 ;
        RECT 75.040 77.800 83.040 77.850 ;
        RECT 74.000 77.620 83.040 77.800 ;
        RECT 74.000 77.600 75.300 77.620 ;
        RECT 74.000 75.300 74.200 77.600 ;
        RECT 74.400 76.700 74.900 77.200 ;
        RECT 84.200 77.100 84.400 79.000 ;
        RECT 85.200 78.580 85.400 80.030 ;
        RECT 86.960 78.920 91.630 79.150 ;
        RECT 91.400 78.900 91.600 78.920 ;
        RECT 92.900 78.580 95.000 78.600 ;
        RECT 85.140 78.400 95.000 78.580 ;
        RECT 85.140 78.350 93.140 78.400 ;
        RECT 93.400 78.090 93.600 78.400 ;
        RECT 94.500 78.100 95.000 78.400 ;
        RECT 93.300 77.900 93.600 78.090 ;
        RECT 93.300 77.550 93.530 77.900 ;
        RECT 85.140 77.200 93.140 77.290 ;
        RECT 84.200 76.800 84.700 77.100 ;
        RECT 82.800 76.710 84.700 76.800 ;
        RECT 74.400 76.350 74.600 76.700 ;
        RECT 75.040 76.600 84.700 76.710 ;
        RECT 84.900 77.060 93.140 77.200 ;
        RECT 84.900 77.000 85.400 77.060 ;
        RECT 75.040 76.480 83.040 76.600 ;
        RECT 84.900 76.400 85.100 77.000 ;
        RECT 74.400 76.100 74.680 76.350 ;
        RECT 74.450 75.550 74.680 76.100 ;
        RECT 83.200 76.200 83.430 76.220 ;
        RECT 84.400 76.200 85.100 76.400 ;
        RECT 95.200 76.200 95.400 81.900 ;
        RECT 83.200 75.700 84.000 76.200 ;
        RECT 83.200 75.680 83.430 75.700 ;
        RECT 75.040 75.300 83.040 75.420 ;
        RECT 74.000 75.190 83.040 75.300 ;
        RECT 74.000 75.100 75.300 75.190 ;
        RECT 74.000 70.500 74.200 75.100 ;
        RECT 74.400 74.300 74.900 74.800 ;
        RECT 84.400 74.300 84.600 76.200 ;
        RECT 91.400 76.150 95.400 76.200 ;
        RECT 86.975 76.000 95.400 76.150 ;
        RECT 86.975 75.920 91.665 76.000 ;
        RECT 95.200 75.600 95.400 76.000 ;
        RECT 92.800 75.580 95.400 75.600 ;
        RECT 85.140 75.400 95.400 75.580 ;
        RECT 85.140 75.350 93.140 75.400 ;
        RECT 93.400 75.090 94.300 75.100 ;
        RECT 93.345 74.600 94.300 75.090 ;
        RECT 93.345 74.550 93.575 74.600 ;
        RECT 74.400 73.920 74.600 74.300 ;
        RECT 82.800 74.280 84.600 74.300 ;
        RECT 75.040 74.100 84.600 74.280 ;
        RECT 75.040 74.050 83.040 74.100 ;
        RECT 74.400 73.120 74.680 73.920 ;
        RECT 83.800 73.800 84.000 74.100 ;
        RECT 85.140 74.060 93.140 74.290 ;
        RECT 83.300 73.790 84.000 73.800 ;
        RECT 83.200 73.300 84.000 73.790 ;
        RECT 83.200 73.250 83.430 73.300 ;
        RECT 85.200 73.150 85.400 74.060 ;
        RECT 86.980 73.700 91.670 73.720 ;
        RECT 95.200 73.700 95.400 75.400 ;
        RECT 86.980 73.500 95.400 73.700 ;
        RECT 86.980 73.490 91.670 73.500 ;
        RECT 74.400 72.900 74.600 73.120 ;
        RECT 75.040 72.900 83.040 72.990 ;
        RECT 85.145 72.920 93.145 73.150 ;
        RECT 74.400 72.760 83.040 72.900 ;
        RECT 74.400 72.700 75.300 72.760 ;
        RECT 93.400 72.660 94.300 72.700 ;
        RECT 74.400 71.800 74.900 72.300 ;
        RECT 93.350 72.200 94.300 72.660 ;
        RECT 84.200 71.900 84.700 72.200 ;
        RECT 93.350 72.120 93.600 72.200 ;
        RECT 82.800 71.850 84.700 71.900 ;
        RECT 74.400 71.490 74.600 71.800 ;
        RECT 75.040 71.700 84.700 71.850 ;
        RECT 75.040 71.620 83.040 71.700 ;
        RECT 74.400 71.300 74.680 71.490 ;
        RECT 74.450 70.690 74.680 71.300 ;
        RECT 83.200 71.300 83.430 71.360 ;
        RECT 83.200 70.820 84.000 71.300 ;
        RECT 83.300 70.800 84.000 70.820 ;
        RECT 75.040 70.500 83.040 70.560 ;
        RECT 74.000 70.330 83.040 70.500 ;
        RECT 74.000 70.300 75.300 70.330 ;
        RECT 74.000 68.100 74.200 70.300 ;
        RECT 74.400 69.400 74.900 69.900 ;
        RECT 84.200 69.500 84.400 71.700 ;
        RECT 85.145 71.630 93.145 71.860 ;
        RECT 85.200 70.170 85.400 71.630 ;
        RECT 86.975 70.510 91.645 70.740 ;
        RECT 93.400 70.200 93.600 72.120 ;
        RECT 92.900 70.170 93.600 70.200 ;
        RECT 85.155 70.000 93.600 70.170 ;
        RECT 85.155 69.940 93.155 70.000 ;
        RECT 94.500 69.700 95.000 69.900 ;
        RECT 93.400 69.680 95.000 69.700 ;
        RECT 82.800 69.420 84.400 69.500 ;
        RECT 74.400 69.060 74.600 69.400 ;
        RECT 75.040 69.300 84.400 69.420 ;
        RECT 75.040 69.190 83.040 69.300 ;
        RECT 74.400 68.900 74.680 69.060 ;
        RECT 74.450 68.260 74.680 68.900 ;
        RECT 83.200 68.900 83.430 68.930 ;
        RECT 83.200 68.400 84.000 68.900 ;
        RECT 84.200 68.800 84.400 69.300 ;
        RECT 93.315 69.400 95.000 69.680 ;
        RECT 93.315 69.140 93.545 69.400 ;
        RECT 85.155 68.800 93.155 68.880 ;
        RECT 84.200 68.650 93.155 68.800 ;
        RECT 84.200 68.600 85.400 68.650 ;
        RECT 83.200 68.390 83.430 68.400 ;
        RECT 75.040 68.100 83.040 68.130 ;
        RECT 74.000 67.900 83.040 68.100 ;
        RECT 74.000 65.600 74.200 67.900 ;
        RECT 74.400 66.900 74.900 67.400 ;
        RECT 84.200 67.000 84.400 68.600 ;
        RECT 95.200 67.800 95.400 73.500 ;
        RECT 91.400 67.750 95.400 67.800 ;
        RECT 86.975 67.600 95.400 67.750 ;
        RECT 86.975 67.520 91.665 67.600 ;
        RECT 95.200 67.200 95.400 67.600 ;
        RECT 92.800 67.180 95.400 67.200 ;
        RECT 82.800 66.990 84.400 67.000 ;
        RECT 74.400 66.630 74.600 66.900 ;
        RECT 75.040 66.800 84.400 66.990 ;
        RECT 85.140 67.000 95.400 67.180 ;
        RECT 85.140 66.950 93.140 67.000 ;
        RECT 75.040 66.760 83.040 66.800 ;
        RECT 74.400 66.400 74.680 66.630 ;
        RECT 74.450 65.830 74.680 66.400 ;
        RECT 83.200 66.000 84.000 66.500 ;
        RECT 83.200 65.960 83.430 66.000 ;
        RECT 75.040 65.600 83.040 65.700 ;
        RECT 74.000 65.470 83.040 65.600 ;
        RECT 74.000 65.400 75.300 65.470 ;
        RECT 74.000 63.200 74.200 65.400 ;
        RECT 74.400 64.500 74.900 65.000 ;
        RECT 84.200 64.600 84.400 66.800 ;
        RECT 93.400 66.690 94.300 66.700 ;
        RECT 93.345 66.200 94.300 66.690 ;
        RECT 93.345 66.150 93.575 66.200 ;
        RECT 85.140 65.660 93.140 65.890 ;
        RECT 85.300 64.780 85.500 65.660 ;
        RECT 95.200 65.400 95.400 67.000 ;
        RECT 91.400 65.350 95.400 65.400 ;
        RECT 86.975 65.200 95.400 65.350 ;
        RECT 86.975 65.120 91.665 65.200 ;
        RECT 82.800 64.560 84.400 64.600 ;
        RECT 74.400 64.200 74.600 64.500 ;
        RECT 75.040 64.400 84.400 64.560 ;
        RECT 85.140 64.550 93.140 64.780 ;
        RECT 75.040 64.330 83.040 64.400 ;
        RECT 93.400 64.290 94.300 64.300 ;
        RECT 74.400 63.900 74.680 64.200 ;
        RECT 83.300 64.070 84.000 64.100 ;
        RECT 74.450 63.400 74.680 63.900 ;
        RECT 83.200 63.600 84.000 64.070 ;
        RECT 93.345 63.800 94.300 64.290 ;
        RECT 93.345 63.750 93.575 63.800 ;
        RECT 83.200 63.530 83.430 63.600 ;
        RECT 85.140 63.400 93.140 63.490 ;
        RECT 75.040 63.200 83.040 63.270 ;
        RECT 74.000 63.040 83.040 63.200 ;
        RECT 84.200 63.260 93.140 63.400 ;
        RECT 84.200 63.200 85.400 63.260 ;
        RECT 74.000 63.000 75.300 63.040 ;
        RECT 74.000 53.700 74.200 63.000 ;
        RECT 74.400 62.500 79.200 62.700 ;
        RECT 74.400 62.100 74.900 62.500 ;
        RECT 76.700 62.100 76.900 62.500 ;
        RECT 74.400 62.080 75.400 62.100 ;
        RECT 76.700 62.080 77.700 62.100 ;
        RECT 74.400 61.900 76.040 62.080 ;
        RECT 74.400 60.195 74.600 61.900 ;
        RECT 75.040 61.850 76.040 61.900 ;
        RECT 76.700 61.900 78.340 62.080 ;
        RECT 76.700 60.195 76.900 61.900 ;
        RECT 77.340 61.850 78.340 61.900 ;
        RECT 79.000 60.195 79.200 62.500 ;
        RECT 80.300 62.080 82.200 62.100 ;
        RECT 79.640 61.900 82.940 62.080 ;
        RECT 79.640 61.850 80.640 61.900 ;
        RECT 81.940 61.850 82.940 61.900 ;
        RECT 74.400 59.900 74.680 60.195 ;
        RECT 76.700 59.900 76.980 60.195 ;
        RECT 79.000 59.900 79.280 60.195 ;
        RECT 74.450 55.445 74.680 59.900 ;
        RECT 76.200 55.800 76.430 59.840 ;
        RECT 75.040 53.700 76.040 53.790 ;
        RECT 74.000 53.560 76.040 53.700 ;
        RECT 74.000 53.500 75.300 53.560 ;
        RECT 75.000 53.300 75.300 53.500 ;
        RECT 75.000 52.800 75.500 53.300 ;
        RECT 76.200 52.600 76.400 55.800 ;
        RECT 76.750 55.445 76.980 59.900 ;
        RECT 78.500 55.800 78.730 59.840 ;
        RECT 77.340 53.560 78.340 53.790 ;
        RECT 77.400 53.300 77.700 53.560 ;
        RECT 77.400 52.800 77.900 53.300 ;
        RECT 78.500 52.600 78.700 55.800 ;
        RECT 79.050 55.700 79.280 59.900 ;
        RECT 80.800 55.800 81.030 59.840 ;
        RECT 79.050 55.445 79.300 55.700 ;
        RECT 79.100 53.300 79.300 55.445 ;
        RECT 79.640 53.560 80.640 53.790 ;
        RECT 79.700 53.300 80.000 53.560 ;
        RECT 79.100 53.100 79.500 53.300 ;
        RECT 76.200 52.100 76.700 52.600 ;
        RECT 78.500 52.100 79.000 52.600 ;
        RECT 79.300 51.900 79.500 53.100 ;
        RECT 79.700 52.800 80.200 53.300 ;
        RECT 80.800 52.600 81.000 55.800 ;
        RECT 80.700 52.100 81.200 52.600 ;
        RECT 81.350 51.900 81.580 58.920 ;
        RECT 79.300 51.700 81.580 51.900 ;
        RECT 80.600 47.500 80.800 51.700 ;
        RECT 81.350 51.620 81.580 51.700 ;
        RECT 83.100 51.975 83.330 58.565 ;
        RECT 83.100 48.700 83.300 51.975 ;
        RECT 84.200 48.700 84.400 63.200 ;
        RECT 95.200 63.000 95.400 65.200 ;
        RECT 91.400 62.950 95.400 63.000 ;
        RECT 86.975 62.800 95.400 62.950 ;
        RECT 86.975 62.720 91.665 62.800 ;
        RECT 95.200 62.400 95.400 62.800 ;
        RECT 92.800 62.380 95.400 62.400 ;
        RECT 85.140 62.200 95.400 62.380 ;
        RECT 85.140 62.150 93.140 62.200 ;
        RECT 93.400 61.890 94.300 61.900 ;
        RECT 93.345 61.400 94.300 61.890 ;
        RECT 93.345 61.350 93.575 61.400 ;
        RECT 85.140 60.860 93.140 61.090 ;
        RECT 85.200 59.985 85.400 60.860 ;
        RECT 95.200 60.600 95.400 62.200 ;
        RECT 91.400 60.555 95.400 60.600 ;
        RECT 86.975 60.400 95.400 60.555 ;
        RECT 86.975 60.325 91.665 60.400 ;
        RECT 85.140 59.755 93.140 59.985 ;
        RECT 93.400 59.495 94.300 59.500 ;
        RECT 93.345 59.000 94.300 59.495 ;
        RECT 93.345 58.955 93.575 59.000 ;
        RECT 85.140 58.600 93.140 58.695 ;
        RECT 94.500 58.600 95.000 58.800 ;
        RECT 85.140 58.465 95.000 58.600 ;
        RECT 92.900 58.400 95.000 58.465 ;
        RECT 94.500 58.300 95.000 58.400 ;
        RECT 95.200 58.100 95.400 60.400 ;
        RECT 88.300 58.050 95.400 58.100 ;
        RECT 88.080 57.900 95.400 58.050 ;
        RECT 88.080 57.820 88.980 57.900 ;
        RECT 85.480 57.500 86.280 57.550 ;
        RECT 82.600 48.690 84.400 48.700 ;
        RECT 81.940 48.500 84.400 48.690 ;
        RECT 84.600 57.320 86.280 57.500 ;
        RECT 88.300 57.480 88.500 57.820 ;
        RECT 89.700 57.550 90.700 57.600 ;
        RECT 84.600 57.300 85.800 57.320 ;
        RECT 84.600 56.900 84.800 57.300 ;
        RECT 88.140 57.250 88.560 57.480 ;
        RECT 89.700 57.400 91.245 57.550 ;
        RECT 85.120 56.900 85.350 56.960 ;
        RECT 84.600 56.700 85.350 56.900 ;
        RECT 81.940 48.460 82.940 48.500 ;
        RECT 82.000 48.200 82.200 48.460 ;
        RECT 82.000 47.700 82.500 48.200 ;
        RECT 84.600 47.500 84.800 56.700 ;
        RECT 85.120 48.960 85.350 56.700 ;
        RECT 86.410 49.300 86.640 56.960 ;
        RECT 88.765 51.500 88.995 55.240 ;
        RECT 88.765 51.200 89.000 51.500 ;
        RECT 86.410 48.960 86.700 49.300 ;
        RECT 88.200 49.190 88.400 49.200 ;
        RECT 88.140 48.960 88.560 49.190 ;
        RECT 85.610 48.570 86.150 48.800 ;
        RECT 85.900 48.300 86.100 48.570 ;
        RECT 85.600 47.800 86.100 48.300 ;
        RECT 86.500 48.300 86.700 48.960 ;
        RECT 86.500 48.000 87.000 48.300 ;
        RECT 88.200 48.000 88.400 48.960 ;
        RECT 86.500 47.800 88.400 48.000 ;
        RECT 80.600 47.300 84.800 47.500 ;
        RECT 85.900 47.600 86.100 47.800 ;
        RECT 88.800 47.600 89.000 51.200 ;
        RECT 85.900 47.400 89.000 47.600 ;
        RECT 89.700 48.700 89.900 57.400 ;
        RECT 90.365 57.320 91.245 57.400 ;
        RECT 93.800 57.000 94.300 57.300 ;
        RECT 90.600 56.980 94.300 57.000 ;
        RECT 90.440 56.800 94.300 56.980 ;
        RECT 94.500 56.800 95.000 57.300 ;
        RECT 90.440 56.750 90.860 56.800 ;
        RECT 94.600 55.100 94.800 56.800 ;
        RECT 91.020 52.700 91.250 54.740 ;
        RECT 91.020 52.500 92.000 52.700 ;
        RECT 91.020 50.700 91.250 52.500 ;
        RECT 91.500 52.200 92.000 52.500 ;
        RECT 93.720 51.400 93.950 55.100 ;
        RECT 93.600 51.100 93.950 51.400 ;
        RECT 94.510 54.800 94.800 55.100 ;
        RECT 94.510 51.100 94.740 54.800 ;
        RECT 95.200 54.265 95.400 57.900 ;
        RECT 95.080 54.000 95.400 54.265 ;
        RECT 95.080 51.575 95.310 54.000 ;
        RECT 89.700 48.690 90.700 48.700 ;
        RECT 89.700 48.500 90.860 48.690 ;
        RECT 84.600 47.200 84.800 47.300 ;
        RECT 89.700 47.200 89.900 48.500 ;
        RECT 90.440 48.460 90.860 48.500 ;
        RECT 84.600 47.000 89.900 47.200 ;
        RECT 93.600 46.800 93.800 51.100 ;
        RECT 94.000 50.665 94.460 50.895 ;
        RECT 94.100 49.900 94.300 50.665 ;
        RECT 94.100 49.200 94.800 49.900 ;
        RECT 94.100 48.200 94.800 48.900 ;
        RECT 73.200 46.600 93.800 46.800 ;
        RECT 43.900 4.600 67.800 4.800 ;
        RECT 73.200 4.800 73.400 46.600 ;
        RECT 86.975 42.500 91.665 42.550 ;
        RECT 97.000 42.500 99.000 84.300 ;
        RECT 74.400 42.000 74.900 42.500 ;
        RECT 86.975 42.320 99.000 42.500 ;
        RECT 91.400 42.300 99.000 42.320 ;
        RECT 82.800 42.000 84.400 42.100 ;
        RECT 95.200 42.000 95.400 42.300 ;
        RECT 74.400 41.640 74.600 42.000 ;
        RECT 75.040 41.900 84.400 42.000 ;
        RECT 92.800 41.980 95.400 42.000 ;
        RECT 75.040 41.770 83.040 41.900 ;
        RECT 74.400 41.500 74.680 41.640 ;
        RECT 74.450 40.840 74.680 41.500 ;
        RECT 83.200 41.500 83.430 41.510 ;
        RECT 83.200 41.000 84.000 41.500 ;
        RECT 83.200 40.970 83.430 41.000 ;
        RECT 75.040 40.600 83.040 40.710 ;
        RECT 74.000 40.480 83.040 40.600 ;
        RECT 74.000 40.400 75.300 40.480 ;
        RECT 74.000 38.200 74.200 40.400 ;
        RECT 74.400 39.500 74.900 40.000 ;
        RECT 84.200 39.600 84.400 41.900 ;
        RECT 85.140 41.800 95.400 41.980 ;
        RECT 85.140 41.750 93.140 41.800 ;
        RECT 93.400 41.490 94.300 41.500 ;
        RECT 93.345 41.000 94.300 41.490 ;
        RECT 93.345 40.950 93.575 41.000 ;
        RECT 85.140 40.460 93.140 40.690 ;
        RECT 82.800 39.570 84.400 39.600 ;
        RECT 74.400 39.210 74.600 39.500 ;
        RECT 75.040 39.400 84.400 39.570 ;
        RECT 85.200 39.550 85.400 40.460 ;
        RECT 86.975 40.100 91.665 40.120 ;
        RECT 95.200 40.100 95.400 41.800 ;
        RECT 86.975 39.900 95.400 40.100 ;
        RECT 86.975 39.890 91.665 39.900 ;
        RECT 75.040 39.340 83.040 39.400 ;
        RECT 74.400 39.000 74.680 39.210 ;
        RECT 83.300 39.080 84.000 39.100 ;
        RECT 74.450 38.410 74.680 39.000 ;
        RECT 83.200 38.600 84.000 39.080 ;
        RECT 83.200 38.540 83.430 38.600 ;
        RECT 75.040 38.200 83.040 38.280 ;
        RECT 74.000 38.050 83.040 38.200 ;
        RECT 74.000 38.000 75.300 38.050 ;
        RECT 74.000 35.800 74.200 38.000 ;
        RECT 74.400 37.100 74.900 37.600 ;
        RECT 84.200 37.200 84.400 39.400 ;
        RECT 85.140 39.320 93.140 39.550 ;
        RECT 93.345 39.000 93.575 39.060 ;
        RECT 93.345 38.520 94.300 39.000 ;
        RECT 93.400 38.500 94.300 38.520 ;
        RECT 85.140 38.030 93.140 38.260 ;
        RECT 82.800 37.140 84.400 37.200 ;
        RECT 74.400 36.780 74.600 37.100 ;
        RECT 75.040 37.000 84.400 37.140 ;
        RECT 75.040 36.910 83.040 37.000 ;
        RECT 74.400 36.600 74.680 36.780 ;
        RECT 83.300 36.650 84.000 36.700 ;
        RECT 74.450 35.980 74.680 36.600 ;
        RECT 83.200 36.200 84.000 36.650 ;
        RECT 83.200 36.110 83.430 36.200 ;
        RECT 75.040 35.800 83.040 35.850 ;
        RECT 74.000 35.620 83.040 35.800 ;
        RECT 74.000 35.600 75.300 35.620 ;
        RECT 74.000 33.300 74.200 35.600 ;
        RECT 74.400 34.700 74.900 35.200 ;
        RECT 84.200 35.100 84.400 37.000 ;
        RECT 85.200 36.580 85.400 38.030 ;
        RECT 86.960 36.920 91.630 37.150 ;
        RECT 91.400 36.900 91.600 36.920 ;
        RECT 92.900 36.580 95.000 36.600 ;
        RECT 85.140 36.400 95.000 36.580 ;
        RECT 85.140 36.350 93.140 36.400 ;
        RECT 93.400 36.090 93.600 36.400 ;
        RECT 94.500 36.100 95.000 36.400 ;
        RECT 93.300 35.900 93.600 36.090 ;
        RECT 93.300 35.550 93.530 35.900 ;
        RECT 85.140 35.200 93.140 35.290 ;
        RECT 84.200 34.800 84.700 35.100 ;
        RECT 82.800 34.710 84.700 34.800 ;
        RECT 74.400 34.350 74.600 34.700 ;
        RECT 75.040 34.600 84.700 34.710 ;
        RECT 84.900 35.060 93.140 35.200 ;
        RECT 84.900 35.000 85.400 35.060 ;
        RECT 75.040 34.480 83.040 34.600 ;
        RECT 84.900 34.400 85.100 35.000 ;
        RECT 74.400 34.100 74.680 34.350 ;
        RECT 74.450 33.550 74.680 34.100 ;
        RECT 83.200 34.200 83.430 34.220 ;
        RECT 84.400 34.200 85.100 34.400 ;
        RECT 95.200 34.200 95.400 39.900 ;
        RECT 83.200 33.700 84.000 34.200 ;
        RECT 83.200 33.680 83.430 33.700 ;
        RECT 75.040 33.300 83.040 33.420 ;
        RECT 74.000 33.190 83.040 33.300 ;
        RECT 74.000 33.100 75.300 33.190 ;
        RECT 74.000 28.500 74.200 33.100 ;
        RECT 74.400 32.300 74.900 32.800 ;
        RECT 84.400 32.300 84.600 34.200 ;
        RECT 91.400 34.150 95.400 34.200 ;
        RECT 86.975 34.000 95.400 34.150 ;
        RECT 86.975 33.920 91.665 34.000 ;
        RECT 95.200 33.600 95.400 34.000 ;
        RECT 92.800 33.580 95.400 33.600 ;
        RECT 85.140 33.400 95.400 33.580 ;
        RECT 85.140 33.350 93.140 33.400 ;
        RECT 93.400 33.090 94.300 33.100 ;
        RECT 93.345 32.600 94.300 33.090 ;
        RECT 93.345 32.550 93.575 32.600 ;
        RECT 74.400 31.920 74.600 32.300 ;
        RECT 82.800 32.280 84.600 32.300 ;
        RECT 75.040 32.100 84.600 32.280 ;
        RECT 75.040 32.050 83.040 32.100 ;
        RECT 74.400 31.120 74.680 31.920 ;
        RECT 83.800 31.800 84.000 32.100 ;
        RECT 85.140 32.060 93.140 32.290 ;
        RECT 83.300 31.790 84.000 31.800 ;
        RECT 83.200 31.300 84.000 31.790 ;
        RECT 83.200 31.250 83.430 31.300 ;
        RECT 85.200 31.150 85.400 32.060 ;
        RECT 86.980 31.700 91.670 31.720 ;
        RECT 95.200 31.700 95.400 33.400 ;
        RECT 86.980 31.500 95.400 31.700 ;
        RECT 86.980 31.490 91.670 31.500 ;
        RECT 74.400 30.900 74.600 31.120 ;
        RECT 75.040 30.900 83.040 30.990 ;
        RECT 85.145 30.920 93.145 31.150 ;
        RECT 74.400 30.760 83.040 30.900 ;
        RECT 74.400 30.700 75.300 30.760 ;
        RECT 93.400 30.660 94.300 30.700 ;
        RECT 74.400 29.800 74.900 30.300 ;
        RECT 93.350 30.200 94.300 30.660 ;
        RECT 84.200 29.900 84.700 30.200 ;
        RECT 93.350 30.120 93.600 30.200 ;
        RECT 82.800 29.850 84.700 29.900 ;
        RECT 74.400 29.490 74.600 29.800 ;
        RECT 75.040 29.700 84.700 29.850 ;
        RECT 75.040 29.620 83.040 29.700 ;
        RECT 74.400 29.300 74.680 29.490 ;
        RECT 74.450 28.690 74.680 29.300 ;
        RECT 83.200 29.300 83.430 29.360 ;
        RECT 83.200 28.820 84.000 29.300 ;
        RECT 83.300 28.800 84.000 28.820 ;
        RECT 75.040 28.500 83.040 28.560 ;
        RECT 74.000 28.330 83.040 28.500 ;
        RECT 74.000 28.300 75.300 28.330 ;
        RECT 74.000 26.100 74.200 28.300 ;
        RECT 74.400 27.400 74.900 27.900 ;
        RECT 84.200 27.500 84.400 29.700 ;
        RECT 85.145 29.630 93.145 29.860 ;
        RECT 85.200 28.170 85.400 29.630 ;
        RECT 86.975 28.510 91.645 28.740 ;
        RECT 93.400 28.200 93.600 30.120 ;
        RECT 92.900 28.170 93.600 28.200 ;
        RECT 85.155 28.000 93.600 28.170 ;
        RECT 85.155 27.940 93.155 28.000 ;
        RECT 94.500 27.700 95.000 27.900 ;
        RECT 93.400 27.680 95.000 27.700 ;
        RECT 82.800 27.420 84.400 27.500 ;
        RECT 74.400 27.060 74.600 27.400 ;
        RECT 75.040 27.300 84.400 27.420 ;
        RECT 75.040 27.190 83.040 27.300 ;
        RECT 74.400 26.900 74.680 27.060 ;
        RECT 74.450 26.260 74.680 26.900 ;
        RECT 83.200 26.900 83.430 26.930 ;
        RECT 83.200 26.400 84.000 26.900 ;
        RECT 84.200 26.800 84.400 27.300 ;
        RECT 93.315 27.400 95.000 27.680 ;
        RECT 93.315 27.140 93.545 27.400 ;
        RECT 85.155 26.800 93.155 26.880 ;
        RECT 84.200 26.650 93.155 26.800 ;
        RECT 84.200 26.600 85.400 26.650 ;
        RECT 83.200 26.390 83.430 26.400 ;
        RECT 75.040 26.100 83.040 26.130 ;
        RECT 74.000 25.900 83.040 26.100 ;
        RECT 74.000 23.600 74.200 25.900 ;
        RECT 74.400 24.900 74.900 25.400 ;
        RECT 84.200 25.000 84.400 26.600 ;
        RECT 95.200 25.800 95.400 31.500 ;
        RECT 91.400 25.750 95.400 25.800 ;
        RECT 86.975 25.600 95.400 25.750 ;
        RECT 86.975 25.520 91.665 25.600 ;
        RECT 95.200 25.200 95.400 25.600 ;
        RECT 92.800 25.180 95.400 25.200 ;
        RECT 82.800 24.990 84.400 25.000 ;
        RECT 74.400 24.630 74.600 24.900 ;
        RECT 75.040 24.800 84.400 24.990 ;
        RECT 85.140 25.000 95.400 25.180 ;
        RECT 85.140 24.950 93.140 25.000 ;
        RECT 75.040 24.760 83.040 24.800 ;
        RECT 74.400 24.400 74.680 24.630 ;
        RECT 74.450 23.830 74.680 24.400 ;
        RECT 83.200 24.000 84.000 24.500 ;
        RECT 83.200 23.960 83.430 24.000 ;
        RECT 75.040 23.600 83.040 23.700 ;
        RECT 74.000 23.470 83.040 23.600 ;
        RECT 74.000 23.400 75.300 23.470 ;
        RECT 74.000 21.200 74.200 23.400 ;
        RECT 74.400 22.500 74.900 23.000 ;
        RECT 84.200 22.600 84.400 24.800 ;
        RECT 93.400 24.690 94.300 24.700 ;
        RECT 93.345 24.200 94.300 24.690 ;
        RECT 93.345 24.150 93.575 24.200 ;
        RECT 85.140 23.660 93.140 23.890 ;
        RECT 85.300 22.780 85.500 23.660 ;
        RECT 95.200 23.400 95.400 25.000 ;
        RECT 91.400 23.350 95.400 23.400 ;
        RECT 86.975 23.200 95.400 23.350 ;
        RECT 86.975 23.120 91.665 23.200 ;
        RECT 82.800 22.560 84.400 22.600 ;
        RECT 74.400 22.200 74.600 22.500 ;
        RECT 75.040 22.400 84.400 22.560 ;
        RECT 85.140 22.550 93.140 22.780 ;
        RECT 75.040 22.330 83.040 22.400 ;
        RECT 93.400 22.290 94.300 22.300 ;
        RECT 74.400 21.900 74.680 22.200 ;
        RECT 83.300 22.070 84.000 22.100 ;
        RECT 74.450 21.400 74.680 21.900 ;
        RECT 83.200 21.600 84.000 22.070 ;
        RECT 93.345 21.800 94.300 22.290 ;
        RECT 93.345 21.750 93.575 21.800 ;
        RECT 83.200 21.530 83.430 21.600 ;
        RECT 85.140 21.400 93.140 21.490 ;
        RECT 75.040 21.200 83.040 21.270 ;
        RECT 74.000 21.040 83.040 21.200 ;
        RECT 84.200 21.260 93.140 21.400 ;
        RECT 84.200 21.200 85.400 21.260 ;
        RECT 74.000 21.000 75.300 21.040 ;
        RECT 74.000 11.700 74.200 21.000 ;
        RECT 74.400 20.500 79.200 20.700 ;
        RECT 74.400 20.100 74.900 20.500 ;
        RECT 76.700 20.100 76.900 20.500 ;
        RECT 74.400 20.080 75.400 20.100 ;
        RECT 76.700 20.080 77.700 20.100 ;
        RECT 74.400 19.900 76.040 20.080 ;
        RECT 74.400 18.195 74.600 19.900 ;
        RECT 75.040 19.850 76.040 19.900 ;
        RECT 76.700 19.900 78.340 20.080 ;
        RECT 76.700 18.195 76.900 19.900 ;
        RECT 77.340 19.850 78.340 19.900 ;
        RECT 79.000 18.195 79.200 20.500 ;
        RECT 80.300 20.080 82.200 20.100 ;
        RECT 79.640 19.900 82.940 20.080 ;
        RECT 79.640 19.850 80.640 19.900 ;
        RECT 81.940 19.850 82.940 19.900 ;
        RECT 74.400 17.900 74.680 18.195 ;
        RECT 76.700 17.900 76.980 18.195 ;
        RECT 79.000 17.900 79.280 18.195 ;
        RECT 74.450 13.445 74.680 17.900 ;
        RECT 76.200 13.800 76.430 17.840 ;
        RECT 75.040 11.700 76.040 11.790 ;
        RECT 74.000 11.560 76.040 11.700 ;
        RECT 74.000 11.500 75.300 11.560 ;
        RECT 75.000 11.300 75.300 11.500 ;
        RECT 75.000 10.800 75.500 11.300 ;
        RECT 76.200 10.600 76.400 13.800 ;
        RECT 76.750 13.445 76.980 17.900 ;
        RECT 78.500 13.800 78.730 17.840 ;
        RECT 77.340 11.560 78.340 11.790 ;
        RECT 77.400 11.300 77.700 11.560 ;
        RECT 77.400 10.800 77.900 11.300 ;
        RECT 78.500 10.600 78.700 13.800 ;
        RECT 79.050 13.700 79.280 17.900 ;
        RECT 80.800 13.800 81.030 17.840 ;
        RECT 79.050 13.445 79.300 13.700 ;
        RECT 79.100 11.300 79.300 13.445 ;
        RECT 79.640 11.560 80.640 11.790 ;
        RECT 79.700 11.300 80.000 11.560 ;
        RECT 79.100 11.100 79.500 11.300 ;
        RECT 76.200 10.100 76.700 10.600 ;
        RECT 78.500 10.100 79.000 10.600 ;
        RECT 79.300 9.900 79.500 11.100 ;
        RECT 79.700 10.800 80.200 11.300 ;
        RECT 80.800 10.600 81.000 13.800 ;
        RECT 80.700 10.100 81.200 10.600 ;
        RECT 81.350 9.900 81.580 16.920 ;
        RECT 79.300 9.700 81.580 9.900 ;
        RECT 80.600 5.500 80.800 9.700 ;
        RECT 81.350 9.620 81.580 9.700 ;
        RECT 83.100 9.975 83.330 16.565 ;
        RECT 83.100 6.700 83.300 9.975 ;
        RECT 84.200 6.700 84.400 21.200 ;
        RECT 95.200 21.000 95.400 23.200 ;
        RECT 91.400 20.950 95.400 21.000 ;
        RECT 86.975 20.800 95.400 20.950 ;
        RECT 86.975 20.720 91.665 20.800 ;
        RECT 95.200 20.400 95.400 20.800 ;
        RECT 92.800 20.380 95.400 20.400 ;
        RECT 85.140 20.200 95.400 20.380 ;
        RECT 85.140 20.150 93.140 20.200 ;
        RECT 93.400 19.890 94.300 19.900 ;
        RECT 93.345 19.400 94.300 19.890 ;
        RECT 93.345 19.350 93.575 19.400 ;
        RECT 85.140 18.860 93.140 19.090 ;
        RECT 85.200 17.985 85.400 18.860 ;
        RECT 95.200 18.600 95.400 20.200 ;
        RECT 91.400 18.555 95.400 18.600 ;
        RECT 86.975 18.400 95.400 18.555 ;
        RECT 86.975 18.325 91.665 18.400 ;
        RECT 85.140 17.755 93.140 17.985 ;
        RECT 93.400 17.495 94.300 17.500 ;
        RECT 93.345 17.000 94.300 17.495 ;
        RECT 93.345 16.955 93.575 17.000 ;
        RECT 85.140 16.600 93.140 16.695 ;
        RECT 94.500 16.600 95.000 16.800 ;
        RECT 85.140 16.465 95.000 16.600 ;
        RECT 92.900 16.400 95.000 16.465 ;
        RECT 94.500 16.300 95.000 16.400 ;
        RECT 95.200 16.100 95.400 18.400 ;
        RECT 88.300 16.050 95.400 16.100 ;
        RECT 88.080 15.900 95.400 16.050 ;
        RECT 88.080 15.820 88.980 15.900 ;
        RECT 85.480 15.500 86.280 15.550 ;
        RECT 82.600 6.690 84.400 6.700 ;
        RECT 81.940 6.500 84.400 6.690 ;
        RECT 84.600 15.320 86.280 15.500 ;
        RECT 88.300 15.480 88.500 15.820 ;
        RECT 89.700 15.550 90.700 15.600 ;
        RECT 84.600 15.300 85.800 15.320 ;
        RECT 84.600 14.900 84.800 15.300 ;
        RECT 88.140 15.250 88.560 15.480 ;
        RECT 89.700 15.400 91.245 15.550 ;
        RECT 85.120 14.900 85.350 14.960 ;
        RECT 84.600 14.700 85.350 14.900 ;
        RECT 81.940 6.460 82.940 6.500 ;
        RECT 82.000 6.200 82.200 6.460 ;
        RECT 82.000 5.700 82.500 6.200 ;
        RECT 84.600 5.500 84.800 14.700 ;
        RECT 85.120 6.960 85.350 14.700 ;
        RECT 86.410 7.300 86.640 14.960 ;
        RECT 88.765 9.500 88.995 13.240 ;
        RECT 88.765 9.200 89.000 9.500 ;
        RECT 86.410 6.960 86.700 7.300 ;
        RECT 88.200 7.190 88.400 7.200 ;
        RECT 88.140 6.960 88.560 7.190 ;
        RECT 85.610 6.570 86.150 6.800 ;
        RECT 85.900 6.300 86.100 6.570 ;
        RECT 85.600 5.800 86.100 6.300 ;
        RECT 86.500 6.300 86.700 6.960 ;
        RECT 86.500 6.000 87.000 6.300 ;
        RECT 88.200 6.000 88.400 6.960 ;
        RECT 86.500 5.800 88.400 6.000 ;
        RECT 80.600 5.300 84.800 5.500 ;
        RECT 85.900 5.600 86.100 5.800 ;
        RECT 88.800 5.600 89.000 9.200 ;
        RECT 85.900 5.400 89.000 5.600 ;
        RECT 89.700 6.700 89.900 15.400 ;
        RECT 90.365 15.320 91.245 15.400 ;
        RECT 93.800 15.000 94.300 15.300 ;
        RECT 90.600 14.980 94.300 15.000 ;
        RECT 90.440 14.800 94.300 14.980 ;
        RECT 94.500 14.800 95.000 15.300 ;
        RECT 90.440 14.750 90.860 14.800 ;
        RECT 94.600 13.100 94.800 14.800 ;
        RECT 91.020 10.700 91.250 12.740 ;
        RECT 91.020 10.500 92.000 10.700 ;
        RECT 91.020 8.700 91.250 10.500 ;
        RECT 91.500 10.200 92.000 10.500 ;
        RECT 93.720 9.400 93.950 13.100 ;
        RECT 93.600 9.100 93.950 9.400 ;
        RECT 94.510 12.800 94.800 13.100 ;
        RECT 94.510 9.100 94.740 12.800 ;
        RECT 95.200 12.265 95.400 15.900 ;
        RECT 95.080 12.000 95.400 12.265 ;
        RECT 95.080 9.575 95.310 12.000 ;
        RECT 89.700 6.690 90.700 6.700 ;
        RECT 89.700 6.500 90.860 6.690 ;
        RECT 84.600 5.200 84.800 5.300 ;
        RECT 89.700 5.200 89.900 6.500 ;
        RECT 90.440 6.460 90.860 6.500 ;
        RECT 84.600 5.000 89.900 5.200 ;
        RECT 93.600 4.800 93.800 9.100 ;
        RECT 94.000 8.665 94.460 8.895 ;
        RECT 94.100 7.900 94.300 8.665 ;
        RECT 94.100 7.200 94.800 7.900 ;
        RECT 94.100 6.200 94.800 6.900 ;
        RECT 97.000 5.000 99.000 42.300 ;
        RECT 73.200 4.600 93.800 4.800 ;
        RECT 43.900 2.000 44.100 4.600 ;
        RECT 73.200 2.000 73.400 4.600 ;
        RECT 43.900 1.800 152.500 2.000 ;
        RECT 151.800 1.300 152.500 1.800 ;
      LAYER met2 ;
        RECT 4.000 210.000 99.000 212.000 ;
        RECT 2.300 207.700 3.000 208.400 ;
        RECT 4.000 187.900 6.000 210.000 ;
        RECT 44.800 209.000 45.500 209.700 ;
        RECT 45.800 209.000 46.500 209.700 ;
        RECT 46.800 209.000 47.500 209.700 ;
        RECT 47.800 209.000 48.500 209.700 ;
        RECT 48.800 209.000 49.500 209.700 ;
        RECT 49.800 209.000 50.500 209.700 ;
        RECT 50.800 209.000 51.500 209.700 ;
        RECT 51.800 209.000 52.500 209.700 ;
        RECT 12.120 207.700 12.620 208.000 ;
        RECT 20.820 207.700 21.320 208.000 ;
        RECT 12.120 207.500 21.320 207.700 ;
        RECT 31.920 207.700 32.420 208.000 ;
        RECT 33.400 207.700 33.900 208.000 ;
        RECT 31.920 207.500 33.920 207.700 ;
        RECT 7.220 207.100 33.920 207.300 ;
        RECT 40.900 207.100 41.600 207.800 ;
        RECT 41.900 207.300 42.600 207.800 ;
        RECT 44.800 207.300 45.000 209.000 ;
        RECT 45.800 208.700 46.000 209.000 ;
        RECT 41.900 207.100 45.000 207.300 ;
        RECT 45.200 208.500 46.000 208.700 ;
        RECT 7.220 206.800 7.720 207.100 ;
        RECT 9.720 206.800 10.220 207.100 ;
        RECT 15.620 206.800 16.120 207.100 ;
        RECT 18.020 206.800 18.520 207.100 ;
        RECT 24.020 206.400 24.520 207.100 ;
        RECT 26.420 206.400 26.920 207.100 ;
        RECT 28.820 206.400 29.320 207.100 ;
        RECT 31.220 206.400 31.720 207.100 ;
        RECT 33.420 206.800 33.920 207.100 ;
        RECT 38.020 204.800 42.920 205.000 ;
        RECT 38.020 204.500 38.520 204.800 ;
        RECT 42.720 200.000 42.920 204.800 ;
        RECT 42.420 199.500 42.920 200.000 ;
        RECT 42.420 198.600 42.920 199.100 ;
        RECT 13.620 197.400 14.120 197.700 ;
        RECT 18.520 197.400 19.020 197.700 ;
        RECT 13.620 197.200 19.020 197.400 ;
        RECT 42.720 197.000 42.920 198.600 ;
        RECT 7.220 196.800 42.920 197.000 ;
        RECT 7.220 196.500 7.720 196.800 ;
        RECT 9.620 196.500 10.120 196.800 ;
        RECT 12.020 196.500 12.520 196.800 ;
        RECT 14.520 196.500 15.020 196.800 ;
        RECT 16.920 196.500 17.420 196.800 ;
        RECT 19.420 196.500 19.920 196.800 ;
        RECT 21.820 196.500 22.320 196.800 ;
        RECT 24.220 196.500 24.720 196.800 ;
        RECT 26.620 196.500 27.120 196.800 ;
        RECT 42.520 195.000 43.020 195.500 ;
        RECT 42.820 194.200 43.020 195.000 ;
        RECT 38.120 194.000 43.020 194.200 ;
        RECT 38.120 193.700 38.620 194.000 ;
        RECT 37.420 192.700 37.920 193.200 ;
        RECT 37.720 190.900 37.920 192.700 ;
        RECT 38.420 192.000 38.620 193.700 ;
        RECT 38.120 191.500 38.620 192.000 ;
        RECT 37.420 190.400 37.920 190.900 ;
        RECT 37.720 188.500 37.920 190.400 ;
        RECT 38.420 189.700 38.620 191.500 ;
        RECT 38.120 189.200 38.620 189.700 ;
        RECT 37.420 188.000 37.920 188.500 ;
        RECT 4.000 187.600 6.720 187.900 ;
        RECT 8.720 187.600 9.220 187.900 ;
        RECT 11.120 187.600 11.620 187.900 ;
        RECT 13.520 187.600 14.020 187.900 ;
        RECT 15.920 187.600 16.420 187.900 ;
        RECT 18.420 187.600 18.920 187.900 ;
        RECT 20.820 187.600 21.320 187.900 ;
        RECT 23.320 187.600 23.820 187.900 ;
        RECT 25.720 187.600 26.220 187.900 ;
        RECT 28.020 187.600 28.520 187.900 ;
        RECT 4.000 187.400 28.520 187.600 ;
        RECT 4.000 187.000 6.000 187.400 ;
        RECT 2.300 181.700 3.000 182.400 ;
        RECT 12.120 181.700 12.620 182.000 ;
        RECT 20.820 181.700 21.320 182.000 ;
        RECT 12.120 181.500 21.320 181.700 ;
        RECT 31.920 181.700 32.420 182.000 ;
        RECT 33.400 181.700 33.900 182.000 ;
        RECT 31.920 181.500 33.920 181.700 ;
        RECT 7.220 181.100 33.920 181.300 ;
        RECT 40.900 181.100 41.600 181.800 ;
        RECT 41.900 181.300 42.600 181.800 ;
        RECT 45.200 181.300 45.400 208.500 ;
        RECT 46.800 208.300 47.000 209.000 ;
        RECT 41.900 181.100 45.400 181.300 ;
        RECT 45.600 208.100 47.000 208.300 ;
        RECT 7.220 180.800 7.720 181.100 ;
        RECT 9.720 180.800 10.220 181.100 ;
        RECT 15.620 180.800 16.120 181.100 ;
        RECT 18.020 180.800 18.520 181.100 ;
        RECT 24.020 180.400 24.520 181.100 ;
        RECT 26.420 180.400 26.920 181.100 ;
        RECT 28.820 180.400 29.320 181.100 ;
        RECT 31.220 180.400 31.720 181.100 ;
        RECT 33.420 180.800 33.920 181.100 ;
        RECT 38.020 178.800 42.920 179.000 ;
        RECT 38.020 178.500 38.520 178.800 ;
        RECT 42.720 174.000 42.920 178.800 ;
        RECT 42.420 173.500 42.920 174.000 ;
        RECT 42.420 172.600 42.920 173.100 ;
        RECT 13.620 171.400 14.120 171.700 ;
        RECT 18.520 171.400 19.020 171.700 ;
        RECT 13.620 171.200 19.020 171.400 ;
        RECT 42.720 171.000 42.920 172.600 ;
        RECT 7.220 170.800 42.920 171.000 ;
        RECT 7.220 170.500 7.720 170.800 ;
        RECT 9.620 170.500 10.120 170.800 ;
        RECT 12.020 170.500 12.520 170.800 ;
        RECT 14.520 170.500 15.020 170.800 ;
        RECT 16.920 170.500 17.420 170.800 ;
        RECT 19.420 170.500 19.920 170.800 ;
        RECT 21.820 170.500 22.320 170.800 ;
        RECT 24.220 170.500 24.720 170.800 ;
        RECT 26.620 170.500 27.120 170.800 ;
        RECT 42.520 169.000 43.020 169.500 ;
        RECT 42.820 168.200 43.020 169.000 ;
        RECT 38.120 168.000 43.020 168.200 ;
        RECT 38.120 167.700 38.620 168.000 ;
        RECT 37.420 166.700 37.920 167.200 ;
        RECT 37.720 164.900 37.920 166.700 ;
        RECT 38.420 166.000 38.620 167.700 ;
        RECT 38.120 165.500 38.620 166.000 ;
        RECT 37.420 164.400 37.920 164.900 ;
        RECT 37.720 162.500 37.920 164.400 ;
        RECT 38.420 163.700 38.620 165.500 ;
        RECT 38.120 163.200 38.620 163.700 ;
        RECT 37.420 162.000 37.920 162.500 ;
        RECT 5.300 161.900 6.000 162.000 ;
        RECT 5.300 161.600 6.720 161.900 ;
        RECT 8.720 161.600 9.220 161.900 ;
        RECT 11.120 161.600 11.620 161.900 ;
        RECT 13.520 161.600 14.020 161.900 ;
        RECT 15.920 161.600 16.420 161.900 ;
        RECT 18.420 161.600 18.920 161.900 ;
        RECT 20.820 161.600 21.320 161.900 ;
        RECT 23.320 161.600 23.820 161.900 ;
        RECT 25.720 161.600 26.220 161.900 ;
        RECT 28.020 161.600 28.520 161.900 ;
        RECT 5.300 161.400 28.520 161.600 ;
        RECT 5.300 161.300 6.000 161.400 ;
        RECT 2.300 155.700 3.000 156.400 ;
        RECT 12.120 155.700 12.620 156.000 ;
        RECT 20.820 155.700 21.320 156.000 ;
        RECT 12.120 155.500 21.320 155.700 ;
        RECT 31.920 155.700 32.420 156.000 ;
        RECT 33.400 155.700 33.900 156.000 ;
        RECT 31.920 155.500 33.920 155.700 ;
        RECT 7.220 155.100 33.920 155.300 ;
        RECT 40.900 155.100 41.600 155.800 ;
        RECT 41.900 155.300 42.600 155.800 ;
        RECT 45.600 155.300 45.800 208.100 ;
        RECT 47.800 207.900 48.000 209.000 ;
        RECT 41.900 155.100 45.800 155.300 ;
        RECT 46.000 207.700 48.000 207.900 ;
        RECT 7.220 154.800 7.720 155.100 ;
        RECT 9.720 154.800 10.220 155.100 ;
        RECT 15.620 154.800 16.120 155.100 ;
        RECT 18.020 154.800 18.520 155.100 ;
        RECT 24.020 154.400 24.520 155.100 ;
        RECT 26.420 154.400 26.920 155.100 ;
        RECT 28.820 154.400 29.320 155.100 ;
        RECT 31.220 154.400 31.720 155.100 ;
        RECT 33.420 154.800 33.920 155.100 ;
        RECT 38.020 152.800 42.920 153.000 ;
        RECT 38.020 152.500 38.520 152.800 ;
        RECT 42.720 148.000 42.920 152.800 ;
        RECT 42.420 147.500 42.920 148.000 ;
        RECT 42.420 146.600 42.920 147.100 ;
        RECT 13.620 145.400 14.120 145.700 ;
        RECT 18.520 145.400 19.020 145.700 ;
        RECT 13.620 145.200 19.020 145.400 ;
        RECT 42.720 145.000 42.920 146.600 ;
        RECT 7.220 144.800 42.920 145.000 ;
        RECT 7.220 144.500 7.720 144.800 ;
        RECT 9.620 144.500 10.120 144.800 ;
        RECT 12.020 144.500 12.520 144.800 ;
        RECT 14.520 144.500 15.020 144.800 ;
        RECT 16.920 144.500 17.420 144.800 ;
        RECT 19.420 144.500 19.920 144.800 ;
        RECT 21.820 144.500 22.320 144.800 ;
        RECT 24.220 144.500 24.720 144.800 ;
        RECT 26.620 144.500 27.120 144.800 ;
        RECT 42.520 143.000 43.020 143.500 ;
        RECT 42.820 142.200 43.020 143.000 ;
        RECT 38.120 142.000 43.020 142.200 ;
        RECT 38.120 141.700 38.620 142.000 ;
        RECT 37.420 140.700 37.920 141.200 ;
        RECT 37.720 138.900 37.920 140.700 ;
        RECT 38.420 140.000 38.620 141.700 ;
        RECT 38.120 139.500 38.620 140.000 ;
        RECT 37.420 138.400 37.920 138.900 ;
        RECT 37.720 136.500 37.920 138.400 ;
        RECT 38.420 137.700 38.620 139.500 ;
        RECT 38.120 137.200 38.620 137.700 ;
        RECT 37.420 136.000 37.920 136.500 ;
        RECT 5.300 135.900 6.000 136.000 ;
        RECT 5.300 135.600 6.720 135.900 ;
        RECT 8.720 135.600 9.220 135.900 ;
        RECT 11.120 135.600 11.620 135.900 ;
        RECT 13.520 135.600 14.020 135.900 ;
        RECT 15.920 135.600 16.420 135.900 ;
        RECT 18.420 135.600 18.920 135.900 ;
        RECT 20.820 135.600 21.320 135.900 ;
        RECT 23.320 135.600 23.820 135.900 ;
        RECT 25.720 135.600 26.220 135.900 ;
        RECT 28.020 135.600 28.520 135.900 ;
        RECT 5.300 135.400 28.520 135.600 ;
        RECT 5.300 135.300 6.000 135.400 ;
        RECT 2.300 129.700 3.000 130.400 ;
        RECT 12.120 129.700 12.620 130.000 ;
        RECT 20.820 129.700 21.320 130.000 ;
        RECT 12.120 129.500 21.320 129.700 ;
        RECT 31.920 129.700 32.420 130.000 ;
        RECT 33.400 129.700 33.900 130.000 ;
        RECT 31.920 129.500 33.920 129.700 ;
        RECT 7.220 129.100 33.920 129.300 ;
        RECT 40.900 129.100 41.600 129.800 ;
        RECT 41.900 129.300 42.600 129.800 ;
        RECT 46.000 129.300 46.200 207.700 ;
        RECT 48.800 207.500 49.000 209.000 ;
        RECT 41.900 129.100 46.200 129.300 ;
        RECT 46.400 207.300 49.000 207.500 ;
        RECT 7.220 128.800 7.720 129.100 ;
        RECT 9.720 128.800 10.220 129.100 ;
        RECT 15.620 128.800 16.120 129.100 ;
        RECT 18.020 128.800 18.520 129.100 ;
        RECT 24.020 128.400 24.520 129.100 ;
        RECT 26.420 128.400 26.920 129.100 ;
        RECT 28.820 128.400 29.320 129.100 ;
        RECT 31.220 128.400 31.720 129.100 ;
        RECT 33.420 128.800 33.920 129.100 ;
        RECT 38.020 126.800 42.920 127.000 ;
        RECT 38.020 126.500 38.520 126.800 ;
        RECT 42.720 122.000 42.920 126.800 ;
        RECT 42.420 121.500 42.920 122.000 ;
        RECT 42.420 120.600 42.920 121.100 ;
        RECT 13.620 119.400 14.120 119.700 ;
        RECT 18.520 119.400 19.020 119.700 ;
        RECT 13.620 119.200 19.020 119.400 ;
        RECT 42.720 119.000 42.920 120.600 ;
        RECT 7.220 118.800 42.920 119.000 ;
        RECT 7.220 118.500 7.720 118.800 ;
        RECT 9.620 118.500 10.120 118.800 ;
        RECT 12.020 118.500 12.520 118.800 ;
        RECT 14.520 118.500 15.020 118.800 ;
        RECT 16.920 118.500 17.420 118.800 ;
        RECT 19.420 118.500 19.920 118.800 ;
        RECT 21.820 118.500 22.320 118.800 ;
        RECT 24.220 118.500 24.720 118.800 ;
        RECT 26.620 118.500 27.120 118.800 ;
        RECT 42.520 117.000 43.020 117.500 ;
        RECT 42.820 116.200 43.020 117.000 ;
        RECT 38.120 116.000 43.020 116.200 ;
        RECT 38.120 115.700 38.620 116.000 ;
        RECT 37.420 114.700 37.920 115.200 ;
        RECT 37.720 112.900 37.920 114.700 ;
        RECT 38.420 114.000 38.620 115.700 ;
        RECT 38.120 113.500 38.620 114.000 ;
        RECT 37.420 112.400 37.920 112.900 ;
        RECT 37.720 110.500 37.920 112.400 ;
        RECT 38.420 111.700 38.620 113.500 ;
        RECT 38.120 111.200 38.620 111.700 ;
        RECT 37.420 110.000 37.920 110.500 ;
        RECT 5.300 109.900 6.000 110.000 ;
        RECT 5.300 109.600 6.720 109.900 ;
        RECT 8.720 109.600 9.220 109.900 ;
        RECT 11.120 109.600 11.620 109.900 ;
        RECT 13.520 109.600 14.020 109.900 ;
        RECT 15.920 109.600 16.420 109.900 ;
        RECT 18.420 109.600 18.920 109.900 ;
        RECT 20.820 109.600 21.320 109.900 ;
        RECT 23.320 109.600 23.820 109.900 ;
        RECT 25.720 109.600 26.220 109.900 ;
        RECT 28.020 109.600 28.520 109.900 ;
        RECT 5.300 109.400 28.520 109.600 ;
        RECT 5.300 109.300 6.000 109.400 ;
        RECT 2.300 103.700 3.000 104.400 ;
        RECT 12.120 103.700 12.620 104.000 ;
        RECT 20.820 103.700 21.320 104.000 ;
        RECT 12.120 103.500 21.320 103.700 ;
        RECT 31.920 103.700 32.420 104.000 ;
        RECT 33.400 103.700 33.900 104.000 ;
        RECT 31.920 103.500 33.920 103.700 ;
        RECT 7.220 103.100 33.920 103.300 ;
        RECT 40.900 103.100 41.600 103.800 ;
        RECT 41.900 103.300 42.600 103.800 ;
        RECT 46.400 103.300 46.600 207.300 ;
        RECT 49.800 207.100 50.000 209.000 ;
        RECT 41.900 103.100 46.600 103.300 ;
        RECT 46.800 206.900 50.000 207.100 ;
        RECT 7.220 102.800 7.720 103.100 ;
        RECT 9.720 102.800 10.220 103.100 ;
        RECT 15.620 102.800 16.120 103.100 ;
        RECT 18.020 102.800 18.520 103.100 ;
        RECT 24.020 102.400 24.520 103.100 ;
        RECT 26.420 102.400 26.920 103.100 ;
        RECT 28.820 102.400 29.320 103.100 ;
        RECT 31.220 102.400 31.720 103.100 ;
        RECT 33.420 102.800 33.920 103.100 ;
        RECT 38.020 100.800 42.920 101.000 ;
        RECT 38.020 100.500 38.520 100.800 ;
        RECT 42.720 96.000 42.920 100.800 ;
        RECT 42.420 95.500 42.920 96.000 ;
        RECT 42.420 94.600 42.920 95.100 ;
        RECT 13.620 93.400 14.120 93.700 ;
        RECT 18.520 93.400 19.020 93.700 ;
        RECT 13.620 93.200 19.020 93.400 ;
        RECT 42.720 93.000 42.920 94.600 ;
        RECT 7.220 92.800 42.920 93.000 ;
        RECT 7.220 92.500 7.720 92.800 ;
        RECT 9.620 92.500 10.120 92.800 ;
        RECT 12.020 92.500 12.520 92.800 ;
        RECT 14.520 92.500 15.020 92.800 ;
        RECT 16.920 92.500 17.420 92.800 ;
        RECT 19.420 92.500 19.920 92.800 ;
        RECT 21.820 92.500 22.320 92.800 ;
        RECT 24.220 92.500 24.720 92.800 ;
        RECT 26.620 92.500 27.120 92.800 ;
        RECT 42.520 91.000 43.020 91.500 ;
        RECT 42.820 90.200 43.020 91.000 ;
        RECT 38.120 90.000 43.020 90.200 ;
        RECT 38.120 89.700 38.620 90.000 ;
        RECT 37.420 88.700 37.920 89.200 ;
        RECT 37.720 86.900 37.920 88.700 ;
        RECT 38.420 88.000 38.620 89.700 ;
        RECT 38.120 87.500 38.620 88.000 ;
        RECT 37.420 86.400 37.920 86.900 ;
        RECT 37.720 84.500 37.920 86.400 ;
        RECT 38.420 85.700 38.620 87.500 ;
        RECT 38.120 85.200 38.620 85.700 ;
        RECT 37.420 84.000 37.920 84.500 ;
        RECT 5.300 83.900 6.000 84.000 ;
        RECT 5.300 83.600 6.720 83.900 ;
        RECT 8.720 83.600 9.220 83.900 ;
        RECT 11.120 83.600 11.620 83.900 ;
        RECT 13.520 83.600 14.020 83.900 ;
        RECT 15.920 83.600 16.420 83.900 ;
        RECT 18.420 83.600 18.920 83.900 ;
        RECT 20.820 83.600 21.320 83.900 ;
        RECT 23.320 83.600 23.820 83.900 ;
        RECT 25.720 83.600 26.220 83.900 ;
        RECT 28.020 83.600 28.520 83.900 ;
        RECT 5.300 83.400 28.520 83.600 ;
        RECT 5.300 83.300 6.000 83.400 ;
        RECT 2.300 77.700 3.000 78.400 ;
        RECT 12.120 77.700 12.620 78.000 ;
        RECT 20.820 77.700 21.320 78.000 ;
        RECT 12.120 77.500 21.320 77.700 ;
        RECT 31.920 77.700 32.420 78.000 ;
        RECT 33.400 77.700 33.900 78.000 ;
        RECT 31.920 77.500 33.920 77.700 ;
        RECT 7.220 77.100 33.920 77.300 ;
        RECT 40.900 77.100 41.600 77.800 ;
        RECT 41.900 77.300 42.600 77.800 ;
        RECT 46.800 77.300 47.000 206.900 ;
        RECT 50.800 206.700 51.000 209.000 ;
        RECT 41.900 77.100 47.000 77.300 ;
        RECT 47.200 206.500 51.000 206.700 ;
        RECT 7.220 76.800 7.720 77.100 ;
        RECT 9.720 76.800 10.220 77.100 ;
        RECT 15.620 76.800 16.120 77.100 ;
        RECT 18.020 76.800 18.520 77.100 ;
        RECT 24.020 76.400 24.520 77.100 ;
        RECT 26.420 76.400 26.920 77.100 ;
        RECT 28.820 76.400 29.320 77.100 ;
        RECT 31.220 76.400 31.720 77.100 ;
        RECT 33.420 76.800 33.920 77.100 ;
        RECT 38.020 74.800 42.920 75.000 ;
        RECT 38.020 74.500 38.520 74.800 ;
        RECT 42.720 70.000 42.920 74.800 ;
        RECT 42.420 69.500 42.920 70.000 ;
        RECT 42.420 68.600 42.920 69.100 ;
        RECT 13.620 67.400 14.120 67.700 ;
        RECT 18.520 67.400 19.020 67.700 ;
        RECT 13.620 67.200 19.020 67.400 ;
        RECT 42.720 67.000 42.920 68.600 ;
        RECT 7.220 66.800 42.920 67.000 ;
        RECT 7.220 66.500 7.720 66.800 ;
        RECT 9.620 66.500 10.120 66.800 ;
        RECT 12.020 66.500 12.520 66.800 ;
        RECT 14.520 66.500 15.020 66.800 ;
        RECT 16.920 66.500 17.420 66.800 ;
        RECT 19.420 66.500 19.920 66.800 ;
        RECT 21.820 66.500 22.320 66.800 ;
        RECT 24.220 66.500 24.720 66.800 ;
        RECT 26.620 66.500 27.120 66.800 ;
        RECT 42.520 65.000 43.020 65.500 ;
        RECT 42.820 64.200 43.020 65.000 ;
        RECT 38.120 64.000 43.020 64.200 ;
        RECT 38.120 63.700 38.620 64.000 ;
        RECT 37.420 62.700 37.920 63.200 ;
        RECT 37.720 60.900 37.920 62.700 ;
        RECT 38.420 62.000 38.620 63.700 ;
        RECT 38.120 61.500 38.620 62.000 ;
        RECT 37.420 60.400 37.920 60.900 ;
        RECT 37.720 58.500 37.920 60.400 ;
        RECT 38.420 59.700 38.620 61.500 ;
        RECT 38.120 59.200 38.620 59.700 ;
        RECT 37.420 58.000 37.920 58.500 ;
        RECT 5.300 57.900 6.000 58.000 ;
        RECT 5.300 57.600 6.720 57.900 ;
        RECT 8.720 57.600 9.220 57.900 ;
        RECT 11.120 57.600 11.620 57.900 ;
        RECT 13.520 57.600 14.020 57.900 ;
        RECT 15.920 57.600 16.420 57.900 ;
        RECT 18.420 57.600 18.920 57.900 ;
        RECT 20.820 57.600 21.320 57.900 ;
        RECT 23.320 57.600 23.820 57.900 ;
        RECT 25.720 57.600 26.220 57.900 ;
        RECT 28.020 57.600 28.520 57.900 ;
        RECT 5.300 57.400 28.520 57.600 ;
        RECT 5.300 57.300 6.000 57.400 ;
        RECT 2.300 51.700 3.000 52.400 ;
        RECT 12.120 51.700 12.620 52.000 ;
        RECT 20.820 51.700 21.320 52.000 ;
        RECT 12.120 51.500 21.320 51.700 ;
        RECT 31.920 51.700 32.420 52.000 ;
        RECT 33.400 51.700 33.900 52.000 ;
        RECT 31.920 51.500 33.920 51.700 ;
        RECT 7.220 51.100 33.920 51.300 ;
        RECT 40.900 51.100 41.600 51.800 ;
        RECT 41.900 51.300 42.600 51.800 ;
        RECT 47.200 51.300 47.400 206.500 ;
        RECT 51.800 206.300 52.000 209.000 ;
        RECT 41.900 51.100 47.400 51.300 ;
        RECT 47.600 206.100 52.000 206.300 ;
        RECT 7.220 50.800 7.720 51.100 ;
        RECT 9.720 50.800 10.220 51.100 ;
        RECT 15.620 50.800 16.120 51.100 ;
        RECT 18.020 50.800 18.520 51.100 ;
        RECT 24.020 50.400 24.520 51.100 ;
        RECT 26.420 50.400 26.920 51.100 ;
        RECT 28.820 50.400 29.320 51.100 ;
        RECT 31.220 50.400 31.720 51.100 ;
        RECT 33.420 50.800 33.920 51.100 ;
        RECT 38.020 48.800 42.920 49.000 ;
        RECT 38.020 48.500 38.520 48.800 ;
        RECT 42.720 44.000 42.920 48.800 ;
        RECT 42.420 43.500 42.920 44.000 ;
        RECT 42.420 42.600 42.920 43.100 ;
        RECT 13.620 41.400 14.120 41.700 ;
        RECT 18.520 41.400 19.020 41.700 ;
        RECT 13.620 41.200 19.020 41.400 ;
        RECT 42.720 41.000 42.920 42.600 ;
        RECT 7.220 40.800 42.920 41.000 ;
        RECT 7.220 40.500 7.720 40.800 ;
        RECT 9.620 40.500 10.120 40.800 ;
        RECT 12.020 40.500 12.520 40.800 ;
        RECT 14.520 40.500 15.020 40.800 ;
        RECT 16.920 40.500 17.420 40.800 ;
        RECT 19.420 40.500 19.920 40.800 ;
        RECT 21.820 40.500 22.320 40.800 ;
        RECT 24.220 40.500 24.720 40.800 ;
        RECT 26.620 40.500 27.120 40.800 ;
        RECT 42.520 39.000 43.020 39.500 ;
        RECT 42.820 38.200 43.020 39.000 ;
        RECT 38.120 38.000 43.020 38.200 ;
        RECT 38.120 37.700 38.620 38.000 ;
        RECT 37.420 36.700 37.920 37.200 ;
        RECT 37.720 34.900 37.920 36.700 ;
        RECT 38.420 36.000 38.620 37.700 ;
        RECT 38.120 35.500 38.620 36.000 ;
        RECT 37.420 34.400 37.920 34.900 ;
        RECT 37.720 32.500 37.920 34.400 ;
        RECT 38.420 33.700 38.620 35.500 ;
        RECT 38.120 33.200 38.620 33.700 ;
        RECT 37.420 32.000 37.920 32.500 ;
        RECT 5.300 31.900 6.000 32.000 ;
        RECT 5.300 31.600 6.720 31.900 ;
        RECT 8.720 31.600 9.220 31.900 ;
        RECT 11.120 31.600 11.620 31.900 ;
        RECT 13.520 31.600 14.020 31.900 ;
        RECT 15.920 31.600 16.420 31.900 ;
        RECT 18.420 31.600 18.920 31.900 ;
        RECT 20.820 31.600 21.320 31.900 ;
        RECT 23.320 31.600 23.820 31.900 ;
        RECT 25.720 31.600 26.220 31.900 ;
        RECT 28.020 31.600 28.520 31.900 ;
        RECT 5.300 31.400 28.520 31.600 ;
        RECT 5.300 31.300 6.000 31.400 ;
        RECT 2.300 25.700 3.000 26.400 ;
        RECT 12.120 25.700 12.620 26.000 ;
        RECT 20.820 25.700 21.320 26.000 ;
        RECT 12.120 25.500 21.320 25.700 ;
        RECT 31.920 25.700 32.420 26.000 ;
        RECT 33.400 25.700 33.900 26.000 ;
        RECT 31.920 25.500 33.920 25.700 ;
        RECT 7.220 25.100 33.920 25.300 ;
        RECT 40.900 25.100 41.600 25.800 ;
        RECT 41.900 25.300 42.600 25.800 ;
        RECT 47.600 25.300 47.800 206.100 ;
        RECT 71.000 168.900 73.000 210.000 ;
        RECT 97.000 168.900 99.000 210.000 ;
        RECT 48.400 168.700 73.000 168.900 ;
        RECT 48.400 168.500 48.600 168.700 ;
        RECT 48.400 168.000 48.900 168.500 ;
        RECT 48.400 166.000 48.600 168.000 ;
        RECT 57.500 167.000 58.000 167.500 ;
        RECT 67.800 167.000 68.300 167.500 ;
        RECT 48.400 165.500 48.900 166.000 ;
        RECT 48.400 163.600 48.600 165.500 ;
        RECT 57.800 165.100 58.000 167.000 ;
        RECT 57.500 164.600 58.000 165.100 ;
        RECT 68.100 165.000 68.300 167.000 ;
        RECT 48.400 163.100 48.900 163.600 ;
        RECT 48.400 161.200 48.600 163.100 ;
        RECT 57.800 162.700 58.000 164.600 ;
        RECT 67.800 164.500 68.300 165.000 ;
        RECT 57.500 162.200 58.000 162.700 ;
        RECT 48.400 160.700 48.900 161.200 ;
        RECT 48.400 158.800 48.600 160.700 ;
        RECT 57.800 160.200 58.000 162.200 ;
        RECT 57.500 159.700 58.000 160.200 ;
        RECT 48.400 158.300 48.900 158.800 ;
        RECT 48.400 156.300 48.600 158.300 ;
        RECT 57.800 157.800 58.000 159.700 ;
        RECT 57.500 157.300 58.000 157.800 ;
        RECT 48.400 155.800 48.900 156.300 ;
        RECT 48.400 153.900 48.600 155.800 ;
        RECT 57.800 155.300 58.000 157.300 ;
        RECT 58.200 160.600 58.700 161.100 ;
        RECT 58.200 156.200 58.400 160.600 ;
        RECT 68.100 159.100 68.300 164.500 ;
        RECT 67.800 158.600 68.300 159.100 ;
        RECT 68.100 156.700 68.300 158.600 ;
        RECT 67.800 156.200 68.300 156.700 ;
        RECT 58.200 155.700 58.700 156.200 ;
        RECT 57.500 154.800 58.000 155.300 ;
        RECT 48.400 153.400 48.900 153.900 ;
        RECT 48.400 151.400 48.600 153.400 ;
        RECT 57.800 152.900 58.000 154.800 ;
        RECT 57.500 152.400 58.000 152.900 ;
        RECT 48.400 150.900 48.900 151.400 ;
        RECT 48.400 149.000 48.600 150.900 ;
        RECT 57.800 150.500 58.000 152.400 ;
        RECT 68.100 150.700 68.300 156.200 ;
        RECT 68.500 162.100 69.000 162.600 ;
        RECT 68.500 153.900 68.700 162.100 ;
        RECT 68.500 153.400 69.000 153.900 ;
        RECT 57.500 150.000 58.000 150.500 ;
        RECT 67.400 150.200 68.300 150.700 ;
        RECT 48.400 148.500 48.900 149.000 ;
        RECT 48.400 146.700 48.600 148.500 ;
        RECT 57.800 148.100 58.000 150.000 ;
        RECT 68.100 148.300 68.300 150.200 ;
        RECT 57.500 147.600 58.000 148.100 ;
        RECT 67.400 147.800 68.300 148.300 ;
        RECT 48.400 146.200 48.900 146.700 ;
        RECT 49.000 137.000 49.500 137.300 ;
        RECT 51.400 137.000 51.900 137.300 ;
        RECT 53.700 137.000 54.200 137.300 ;
        RECT 49.000 136.800 54.200 137.000 ;
        RECT 50.200 136.300 50.700 136.600 ;
        RECT 52.500 136.300 53.000 136.600 ;
        RECT 54.700 136.300 55.200 136.600 ;
        RECT 50.200 136.100 55.200 136.300 ;
        RECT 55.000 131.900 55.200 136.100 ;
        RECT 56.000 131.900 56.500 132.200 ;
        RECT 55.000 131.700 56.500 131.900 ;
        RECT 57.800 132.000 58.000 147.600 ;
        RECT 68.100 145.900 68.300 147.800 ;
        RECT 67.400 145.400 68.300 145.900 ;
        RECT 68.100 143.500 68.300 145.400 ;
        RECT 67.400 143.000 68.300 143.500 ;
        RECT 68.100 141.300 68.300 143.000 ;
        RECT 67.800 140.800 68.300 141.300 ;
        RECT 68.500 142.300 69.000 142.800 ;
        RECT 68.500 141.300 68.700 142.300 ;
        RECT 68.500 140.800 69.000 141.300 ;
        RECT 65.500 136.200 66.000 136.700 ;
        RECT 59.600 132.000 60.100 132.300 ;
        RECT 57.800 131.800 60.100 132.000 ;
        RECT 60.500 132.000 61.000 132.300 ;
        RECT 65.800 132.000 66.000 136.200 ;
        RECT 68.100 133.200 68.800 133.900 ;
        RECT 68.100 132.200 68.800 132.900 ;
        RECT 60.500 131.800 66.000 132.000 ;
        RECT 71.000 126.900 73.000 168.700 ;
        RECT 74.400 168.700 99.000 168.900 ;
        RECT 74.400 168.500 74.600 168.700 ;
        RECT 74.400 168.000 74.900 168.500 ;
        RECT 74.400 166.000 74.600 168.000 ;
        RECT 83.500 167.000 84.000 167.500 ;
        RECT 93.800 167.000 94.300 167.500 ;
        RECT 74.400 165.500 74.900 166.000 ;
        RECT 74.400 163.600 74.600 165.500 ;
        RECT 83.800 165.100 84.000 167.000 ;
        RECT 83.500 164.600 84.000 165.100 ;
        RECT 94.100 165.000 94.300 167.000 ;
        RECT 74.400 163.100 74.900 163.600 ;
        RECT 74.400 161.200 74.600 163.100 ;
        RECT 83.800 162.700 84.000 164.600 ;
        RECT 93.800 164.500 94.300 165.000 ;
        RECT 83.500 162.200 84.000 162.700 ;
        RECT 74.400 160.700 74.900 161.200 ;
        RECT 74.400 158.800 74.600 160.700 ;
        RECT 83.800 160.200 84.000 162.200 ;
        RECT 83.500 159.700 84.000 160.200 ;
        RECT 74.400 158.300 74.900 158.800 ;
        RECT 74.400 156.300 74.600 158.300 ;
        RECT 83.800 157.800 84.000 159.700 ;
        RECT 83.500 157.300 84.000 157.800 ;
        RECT 74.400 155.800 74.900 156.300 ;
        RECT 74.400 153.900 74.600 155.800 ;
        RECT 83.800 155.300 84.000 157.300 ;
        RECT 84.200 160.600 84.700 161.100 ;
        RECT 84.200 156.200 84.400 160.600 ;
        RECT 94.100 159.100 94.300 164.500 ;
        RECT 93.800 158.600 94.300 159.100 ;
        RECT 94.100 156.700 94.300 158.600 ;
        RECT 93.800 156.200 94.300 156.700 ;
        RECT 84.200 155.700 84.700 156.200 ;
        RECT 83.500 154.800 84.000 155.300 ;
        RECT 74.400 153.400 74.900 153.900 ;
        RECT 74.400 151.400 74.600 153.400 ;
        RECT 83.800 152.900 84.000 154.800 ;
        RECT 83.500 152.400 84.000 152.900 ;
        RECT 74.400 150.900 74.900 151.400 ;
        RECT 74.400 149.000 74.600 150.900 ;
        RECT 83.800 150.500 84.000 152.400 ;
        RECT 94.100 150.700 94.300 156.200 ;
        RECT 94.500 162.100 95.000 162.600 ;
        RECT 94.500 153.900 94.700 162.100 ;
        RECT 94.500 153.400 95.000 153.900 ;
        RECT 83.500 150.000 84.000 150.500 ;
        RECT 93.400 150.200 94.300 150.700 ;
        RECT 74.400 148.500 74.900 149.000 ;
        RECT 74.400 146.700 74.600 148.500 ;
        RECT 83.800 148.100 84.000 150.000 ;
        RECT 94.100 148.300 94.300 150.200 ;
        RECT 83.500 147.600 84.000 148.100 ;
        RECT 93.400 147.800 94.300 148.300 ;
        RECT 74.400 146.200 74.900 146.700 ;
        RECT 75.000 137.000 75.500 137.300 ;
        RECT 77.400 137.000 77.900 137.300 ;
        RECT 79.700 137.000 80.200 137.300 ;
        RECT 75.000 136.800 80.200 137.000 ;
        RECT 76.200 136.300 76.700 136.600 ;
        RECT 78.500 136.300 79.000 136.600 ;
        RECT 80.700 136.300 81.200 136.600 ;
        RECT 76.200 136.100 81.200 136.300 ;
        RECT 81.000 131.900 81.200 136.100 ;
        RECT 82.000 131.900 82.500 132.200 ;
        RECT 81.000 131.700 82.500 131.900 ;
        RECT 83.800 132.000 84.000 147.600 ;
        RECT 94.100 145.900 94.300 147.800 ;
        RECT 93.400 145.400 94.300 145.900 ;
        RECT 94.100 143.500 94.300 145.400 ;
        RECT 93.400 143.000 94.300 143.500 ;
        RECT 94.100 141.300 94.300 143.000 ;
        RECT 93.800 140.800 94.300 141.300 ;
        RECT 94.500 142.300 95.000 142.800 ;
        RECT 94.500 141.300 94.700 142.300 ;
        RECT 94.500 140.800 95.000 141.300 ;
        RECT 91.500 136.200 92.000 136.700 ;
        RECT 85.600 132.000 86.100 132.300 ;
        RECT 83.800 131.800 86.100 132.000 ;
        RECT 86.500 132.000 87.000 132.300 ;
        RECT 91.800 132.000 92.000 136.200 ;
        RECT 94.100 133.200 94.800 133.900 ;
        RECT 94.100 132.200 94.800 132.900 ;
        RECT 86.500 131.800 92.000 132.000 ;
        RECT 97.000 126.900 99.000 168.700 ;
        RECT 48.400 126.700 73.000 126.900 ;
        RECT 48.400 126.500 48.600 126.700 ;
        RECT 48.400 126.000 48.900 126.500 ;
        RECT 48.400 124.000 48.600 126.000 ;
        RECT 57.500 125.000 58.000 125.500 ;
        RECT 67.800 125.000 68.300 125.500 ;
        RECT 48.400 123.500 48.900 124.000 ;
        RECT 48.400 121.600 48.600 123.500 ;
        RECT 57.800 123.100 58.000 125.000 ;
        RECT 57.500 122.600 58.000 123.100 ;
        RECT 68.100 123.000 68.300 125.000 ;
        RECT 48.400 121.100 48.900 121.600 ;
        RECT 48.400 119.200 48.600 121.100 ;
        RECT 57.800 120.700 58.000 122.600 ;
        RECT 67.800 122.500 68.300 123.000 ;
        RECT 57.500 120.200 58.000 120.700 ;
        RECT 48.400 118.700 48.900 119.200 ;
        RECT 48.400 116.800 48.600 118.700 ;
        RECT 57.800 118.200 58.000 120.200 ;
        RECT 57.500 117.700 58.000 118.200 ;
        RECT 48.400 116.300 48.900 116.800 ;
        RECT 48.400 114.300 48.600 116.300 ;
        RECT 57.800 115.800 58.000 117.700 ;
        RECT 57.500 115.300 58.000 115.800 ;
        RECT 48.400 113.800 48.900 114.300 ;
        RECT 48.400 111.900 48.600 113.800 ;
        RECT 57.800 113.300 58.000 115.300 ;
        RECT 58.200 118.600 58.700 119.100 ;
        RECT 58.200 114.200 58.400 118.600 ;
        RECT 68.100 117.100 68.300 122.500 ;
        RECT 67.800 116.600 68.300 117.100 ;
        RECT 68.100 114.700 68.300 116.600 ;
        RECT 67.800 114.200 68.300 114.700 ;
        RECT 58.200 113.700 58.700 114.200 ;
        RECT 57.500 112.800 58.000 113.300 ;
        RECT 48.400 111.400 48.900 111.900 ;
        RECT 48.400 109.400 48.600 111.400 ;
        RECT 57.800 110.900 58.000 112.800 ;
        RECT 57.500 110.400 58.000 110.900 ;
        RECT 48.400 108.900 48.900 109.400 ;
        RECT 48.400 107.000 48.600 108.900 ;
        RECT 57.800 108.500 58.000 110.400 ;
        RECT 68.100 108.700 68.300 114.200 ;
        RECT 68.500 120.100 69.000 120.600 ;
        RECT 68.500 111.900 68.700 120.100 ;
        RECT 68.500 111.400 69.000 111.900 ;
        RECT 57.500 108.000 58.000 108.500 ;
        RECT 67.400 108.200 68.300 108.700 ;
        RECT 48.400 106.500 48.900 107.000 ;
        RECT 48.400 104.700 48.600 106.500 ;
        RECT 57.800 106.100 58.000 108.000 ;
        RECT 68.100 106.300 68.300 108.200 ;
        RECT 57.500 105.600 58.000 106.100 ;
        RECT 67.400 105.800 68.300 106.300 ;
        RECT 48.400 104.200 48.900 104.700 ;
        RECT 49.000 95.000 49.500 95.300 ;
        RECT 51.400 95.000 51.900 95.300 ;
        RECT 53.700 95.000 54.200 95.300 ;
        RECT 49.000 94.800 54.200 95.000 ;
        RECT 50.200 94.300 50.700 94.600 ;
        RECT 52.500 94.300 53.000 94.600 ;
        RECT 54.700 94.300 55.200 94.600 ;
        RECT 50.200 94.100 55.200 94.300 ;
        RECT 55.000 89.900 55.200 94.100 ;
        RECT 56.000 89.900 56.500 90.200 ;
        RECT 55.000 89.700 56.500 89.900 ;
        RECT 57.800 90.000 58.000 105.600 ;
        RECT 68.100 103.900 68.300 105.800 ;
        RECT 67.400 103.400 68.300 103.900 ;
        RECT 68.100 101.500 68.300 103.400 ;
        RECT 67.400 101.000 68.300 101.500 ;
        RECT 68.100 99.300 68.300 101.000 ;
        RECT 67.800 98.800 68.300 99.300 ;
        RECT 68.500 100.300 69.000 100.800 ;
        RECT 68.500 99.300 68.700 100.300 ;
        RECT 68.500 98.800 69.000 99.300 ;
        RECT 65.500 94.200 66.000 94.700 ;
        RECT 59.600 90.000 60.100 90.300 ;
        RECT 57.800 89.800 60.100 90.000 ;
        RECT 60.500 90.000 61.000 90.300 ;
        RECT 65.800 90.000 66.000 94.200 ;
        RECT 68.100 91.200 68.800 91.900 ;
        RECT 68.100 90.200 68.800 90.900 ;
        RECT 60.500 89.800 66.000 90.000 ;
        RECT 71.000 84.900 73.000 126.700 ;
        RECT 74.400 126.700 99.000 126.900 ;
        RECT 74.400 126.500 74.600 126.700 ;
        RECT 74.400 126.000 74.900 126.500 ;
        RECT 74.400 124.000 74.600 126.000 ;
        RECT 83.500 125.000 84.000 125.500 ;
        RECT 93.800 125.000 94.300 125.500 ;
        RECT 74.400 123.500 74.900 124.000 ;
        RECT 74.400 121.600 74.600 123.500 ;
        RECT 83.800 123.100 84.000 125.000 ;
        RECT 83.500 122.600 84.000 123.100 ;
        RECT 94.100 123.000 94.300 125.000 ;
        RECT 74.400 121.100 74.900 121.600 ;
        RECT 74.400 119.200 74.600 121.100 ;
        RECT 83.800 120.700 84.000 122.600 ;
        RECT 93.800 122.500 94.300 123.000 ;
        RECT 83.500 120.200 84.000 120.700 ;
        RECT 74.400 118.700 74.900 119.200 ;
        RECT 74.400 116.800 74.600 118.700 ;
        RECT 83.800 118.200 84.000 120.200 ;
        RECT 83.500 117.700 84.000 118.200 ;
        RECT 74.400 116.300 74.900 116.800 ;
        RECT 74.400 114.300 74.600 116.300 ;
        RECT 83.800 115.800 84.000 117.700 ;
        RECT 83.500 115.300 84.000 115.800 ;
        RECT 74.400 113.800 74.900 114.300 ;
        RECT 74.400 111.900 74.600 113.800 ;
        RECT 83.800 113.300 84.000 115.300 ;
        RECT 84.200 118.600 84.700 119.100 ;
        RECT 84.200 114.200 84.400 118.600 ;
        RECT 94.100 117.100 94.300 122.500 ;
        RECT 93.800 116.600 94.300 117.100 ;
        RECT 94.100 114.700 94.300 116.600 ;
        RECT 93.800 114.200 94.300 114.700 ;
        RECT 84.200 113.700 84.700 114.200 ;
        RECT 83.500 112.800 84.000 113.300 ;
        RECT 74.400 111.400 74.900 111.900 ;
        RECT 74.400 109.400 74.600 111.400 ;
        RECT 83.800 110.900 84.000 112.800 ;
        RECT 83.500 110.400 84.000 110.900 ;
        RECT 74.400 108.900 74.900 109.400 ;
        RECT 74.400 107.000 74.600 108.900 ;
        RECT 83.800 108.500 84.000 110.400 ;
        RECT 94.100 108.700 94.300 114.200 ;
        RECT 94.500 120.100 95.000 120.600 ;
        RECT 94.500 111.900 94.700 120.100 ;
        RECT 94.500 111.400 95.000 111.900 ;
        RECT 83.500 108.000 84.000 108.500 ;
        RECT 93.400 108.200 94.300 108.700 ;
        RECT 74.400 106.500 74.900 107.000 ;
        RECT 74.400 104.700 74.600 106.500 ;
        RECT 83.800 106.100 84.000 108.000 ;
        RECT 94.100 106.300 94.300 108.200 ;
        RECT 83.500 105.600 84.000 106.100 ;
        RECT 93.400 105.800 94.300 106.300 ;
        RECT 74.400 104.200 74.900 104.700 ;
        RECT 75.000 95.000 75.500 95.300 ;
        RECT 77.400 95.000 77.900 95.300 ;
        RECT 79.700 95.000 80.200 95.300 ;
        RECT 75.000 94.800 80.200 95.000 ;
        RECT 76.200 94.300 76.700 94.600 ;
        RECT 78.500 94.300 79.000 94.600 ;
        RECT 80.700 94.300 81.200 94.600 ;
        RECT 76.200 94.100 81.200 94.300 ;
        RECT 81.000 89.900 81.200 94.100 ;
        RECT 82.000 89.900 82.500 90.200 ;
        RECT 81.000 89.700 82.500 89.900 ;
        RECT 83.800 90.000 84.000 105.600 ;
        RECT 94.100 103.900 94.300 105.800 ;
        RECT 93.400 103.400 94.300 103.900 ;
        RECT 94.100 101.500 94.300 103.400 ;
        RECT 93.400 101.000 94.300 101.500 ;
        RECT 94.100 99.300 94.300 101.000 ;
        RECT 93.800 98.800 94.300 99.300 ;
        RECT 94.500 100.300 95.000 100.800 ;
        RECT 94.500 99.300 94.700 100.300 ;
        RECT 94.500 98.800 95.000 99.300 ;
        RECT 91.500 94.200 92.000 94.700 ;
        RECT 85.600 90.000 86.100 90.300 ;
        RECT 83.800 89.800 86.100 90.000 ;
        RECT 86.500 90.000 87.000 90.300 ;
        RECT 91.800 90.000 92.000 94.200 ;
        RECT 94.100 91.200 94.800 91.900 ;
        RECT 94.100 90.200 94.800 90.900 ;
        RECT 86.500 89.800 92.000 90.000 ;
        RECT 97.000 84.900 99.000 126.700 ;
        RECT 48.400 84.700 73.000 84.900 ;
        RECT 48.400 84.500 48.600 84.700 ;
        RECT 48.400 84.000 48.900 84.500 ;
        RECT 48.400 82.000 48.600 84.000 ;
        RECT 57.500 83.000 58.000 83.500 ;
        RECT 67.800 83.000 68.300 83.500 ;
        RECT 48.400 81.500 48.900 82.000 ;
        RECT 48.400 79.600 48.600 81.500 ;
        RECT 57.800 81.100 58.000 83.000 ;
        RECT 57.500 80.600 58.000 81.100 ;
        RECT 68.100 81.000 68.300 83.000 ;
        RECT 48.400 79.100 48.900 79.600 ;
        RECT 48.400 77.200 48.600 79.100 ;
        RECT 57.800 78.700 58.000 80.600 ;
        RECT 67.800 80.500 68.300 81.000 ;
        RECT 57.500 78.200 58.000 78.700 ;
        RECT 48.400 76.700 48.900 77.200 ;
        RECT 48.400 74.800 48.600 76.700 ;
        RECT 57.800 76.200 58.000 78.200 ;
        RECT 57.500 75.700 58.000 76.200 ;
        RECT 48.400 74.300 48.900 74.800 ;
        RECT 48.400 72.300 48.600 74.300 ;
        RECT 57.800 73.800 58.000 75.700 ;
        RECT 57.500 73.300 58.000 73.800 ;
        RECT 48.400 71.800 48.900 72.300 ;
        RECT 48.400 69.900 48.600 71.800 ;
        RECT 57.800 71.300 58.000 73.300 ;
        RECT 58.200 76.600 58.700 77.100 ;
        RECT 58.200 72.200 58.400 76.600 ;
        RECT 68.100 75.100 68.300 80.500 ;
        RECT 67.800 74.600 68.300 75.100 ;
        RECT 68.100 72.700 68.300 74.600 ;
        RECT 67.800 72.200 68.300 72.700 ;
        RECT 58.200 71.700 58.700 72.200 ;
        RECT 57.500 70.800 58.000 71.300 ;
        RECT 48.400 69.400 48.900 69.900 ;
        RECT 48.400 67.400 48.600 69.400 ;
        RECT 57.800 68.900 58.000 70.800 ;
        RECT 57.500 68.400 58.000 68.900 ;
        RECT 48.400 66.900 48.900 67.400 ;
        RECT 48.400 65.000 48.600 66.900 ;
        RECT 57.800 66.500 58.000 68.400 ;
        RECT 68.100 66.700 68.300 72.200 ;
        RECT 68.500 78.100 69.000 78.600 ;
        RECT 68.500 69.900 68.700 78.100 ;
        RECT 68.500 69.400 69.000 69.900 ;
        RECT 57.500 66.000 58.000 66.500 ;
        RECT 67.400 66.200 68.300 66.700 ;
        RECT 48.400 64.500 48.900 65.000 ;
        RECT 48.400 62.700 48.600 64.500 ;
        RECT 57.800 64.100 58.000 66.000 ;
        RECT 68.100 64.300 68.300 66.200 ;
        RECT 57.500 63.600 58.000 64.100 ;
        RECT 67.400 63.800 68.300 64.300 ;
        RECT 48.400 62.200 48.900 62.700 ;
        RECT 49.000 53.000 49.500 53.300 ;
        RECT 51.400 53.000 51.900 53.300 ;
        RECT 53.700 53.000 54.200 53.300 ;
        RECT 49.000 52.800 54.200 53.000 ;
        RECT 50.200 52.300 50.700 52.600 ;
        RECT 52.500 52.300 53.000 52.600 ;
        RECT 54.700 52.300 55.200 52.600 ;
        RECT 50.200 52.100 55.200 52.300 ;
        RECT 55.000 47.900 55.200 52.100 ;
        RECT 56.000 47.900 56.500 48.200 ;
        RECT 55.000 47.700 56.500 47.900 ;
        RECT 57.800 48.000 58.000 63.600 ;
        RECT 68.100 61.900 68.300 63.800 ;
        RECT 67.400 61.400 68.300 61.900 ;
        RECT 68.100 59.500 68.300 61.400 ;
        RECT 67.400 59.000 68.300 59.500 ;
        RECT 68.100 57.300 68.300 59.000 ;
        RECT 67.800 56.800 68.300 57.300 ;
        RECT 68.500 58.300 69.000 58.800 ;
        RECT 68.500 57.300 68.700 58.300 ;
        RECT 68.500 56.800 69.000 57.300 ;
        RECT 65.500 52.200 66.000 52.700 ;
        RECT 59.600 48.000 60.100 48.300 ;
        RECT 57.800 47.800 60.100 48.000 ;
        RECT 60.500 48.000 61.000 48.300 ;
        RECT 65.800 48.000 66.000 52.200 ;
        RECT 68.100 49.200 68.800 49.900 ;
        RECT 68.100 48.200 68.800 48.900 ;
        RECT 60.500 47.800 66.000 48.000 ;
        RECT 71.000 42.900 73.000 84.700 ;
        RECT 74.400 84.700 99.000 84.900 ;
        RECT 74.400 84.500 74.600 84.700 ;
        RECT 74.400 84.000 74.900 84.500 ;
        RECT 74.400 82.000 74.600 84.000 ;
        RECT 83.500 83.000 84.000 83.500 ;
        RECT 93.800 83.000 94.300 83.500 ;
        RECT 74.400 81.500 74.900 82.000 ;
        RECT 74.400 79.600 74.600 81.500 ;
        RECT 83.800 81.100 84.000 83.000 ;
        RECT 83.500 80.600 84.000 81.100 ;
        RECT 94.100 81.000 94.300 83.000 ;
        RECT 74.400 79.100 74.900 79.600 ;
        RECT 74.400 77.200 74.600 79.100 ;
        RECT 83.800 78.700 84.000 80.600 ;
        RECT 93.800 80.500 94.300 81.000 ;
        RECT 83.500 78.200 84.000 78.700 ;
        RECT 74.400 76.700 74.900 77.200 ;
        RECT 74.400 74.800 74.600 76.700 ;
        RECT 83.800 76.200 84.000 78.200 ;
        RECT 83.500 75.700 84.000 76.200 ;
        RECT 74.400 74.300 74.900 74.800 ;
        RECT 74.400 72.300 74.600 74.300 ;
        RECT 83.800 73.800 84.000 75.700 ;
        RECT 83.500 73.300 84.000 73.800 ;
        RECT 74.400 71.800 74.900 72.300 ;
        RECT 74.400 69.900 74.600 71.800 ;
        RECT 83.800 71.300 84.000 73.300 ;
        RECT 84.200 76.600 84.700 77.100 ;
        RECT 84.200 72.200 84.400 76.600 ;
        RECT 94.100 75.100 94.300 80.500 ;
        RECT 93.800 74.600 94.300 75.100 ;
        RECT 94.100 72.700 94.300 74.600 ;
        RECT 93.800 72.200 94.300 72.700 ;
        RECT 84.200 71.700 84.700 72.200 ;
        RECT 83.500 70.800 84.000 71.300 ;
        RECT 74.400 69.400 74.900 69.900 ;
        RECT 74.400 67.400 74.600 69.400 ;
        RECT 83.800 68.900 84.000 70.800 ;
        RECT 83.500 68.400 84.000 68.900 ;
        RECT 74.400 66.900 74.900 67.400 ;
        RECT 74.400 65.000 74.600 66.900 ;
        RECT 83.800 66.500 84.000 68.400 ;
        RECT 94.100 66.700 94.300 72.200 ;
        RECT 94.500 78.100 95.000 78.600 ;
        RECT 94.500 69.900 94.700 78.100 ;
        RECT 94.500 69.400 95.000 69.900 ;
        RECT 83.500 66.000 84.000 66.500 ;
        RECT 93.400 66.200 94.300 66.700 ;
        RECT 74.400 64.500 74.900 65.000 ;
        RECT 74.400 62.700 74.600 64.500 ;
        RECT 83.800 64.100 84.000 66.000 ;
        RECT 94.100 64.300 94.300 66.200 ;
        RECT 83.500 63.600 84.000 64.100 ;
        RECT 93.400 63.800 94.300 64.300 ;
        RECT 74.400 62.200 74.900 62.700 ;
        RECT 75.000 53.000 75.500 53.300 ;
        RECT 77.400 53.000 77.900 53.300 ;
        RECT 79.700 53.000 80.200 53.300 ;
        RECT 75.000 52.800 80.200 53.000 ;
        RECT 76.200 52.300 76.700 52.600 ;
        RECT 78.500 52.300 79.000 52.600 ;
        RECT 80.700 52.300 81.200 52.600 ;
        RECT 76.200 52.100 81.200 52.300 ;
        RECT 81.000 47.900 81.200 52.100 ;
        RECT 82.000 47.900 82.500 48.200 ;
        RECT 81.000 47.700 82.500 47.900 ;
        RECT 83.800 48.000 84.000 63.600 ;
        RECT 94.100 61.900 94.300 63.800 ;
        RECT 93.400 61.400 94.300 61.900 ;
        RECT 94.100 59.500 94.300 61.400 ;
        RECT 93.400 59.000 94.300 59.500 ;
        RECT 94.100 57.300 94.300 59.000 ;
        RECT 93.800 56.800 94.300 57.300 ;
        RECT 94.500 58.300 95.000 58.800 ;
        RECT 94.500 57.300 94.700 58.300 ;
        RECT 94.500 56.800 95.000 57.300 ;
        RECT 91.500 52.200 92.000 52.700 ;
        RECT 85.600 48.000 86.100 48.300 ;
        RECT 83.800 47.800 86.100 48.000 ;
        RECT 86.500 48.000 87.000 48.300 ;
        RECT 91.800 48.000 92.000 52.200 ;
        RECT 94.100 49.200 94.800 49.900 ;
        RECT 94.100 48.200 94.800 48.900 ;
        RECT 86.500 47.800 92.000 48.000 ;
        RECT 97.000 42.900 99.000 84.700 ;
        RECT 41.900 25.100 47.800 25.300 ;
        RECT 48.400 42.700 73.000 42.900 ;
        RECT 48.400 42.500 48.600 42.700 ;
        RECT 48.400 42.000 48.900 42.500 ;
        RECT 48.400 40.000 48.600 42.000 ;
        RECT 57.500 41.000 58.000 41.500 ;
        RECT 67.800 41.000 68.300 41.500 ;
        RECT 48.400 39.500 48.900 40.000 ;
        RECT 48.400 37.600 48.600 39.500 ;
        RECT 57.800 39.100 58.000 41.000 ;
        RECT 57.500 38.600 58.000 39.100 ;
        RECT 68.100 39.000 68.300 41.000 ;
        RECT 48.400 37.100 48.900 37.600 ;
        RECT 48.400 35.200 48.600 37.100 ;
        RECT 57.800 36.700 58.000 38.600 ;
        RECT 67.800 38.500 68.300 39.000 ;
        RECT 57.500 36.200 58.000 36.700 ;
        RECT 48.400 34.700 48.900 35.200 ;
        RECT 48.400 32.800 48.600 34.700 ;
        RECT 57.800 34.200 58.000 36.200 ;
        RECT 57.500 33.700 58.000 34.200 ;
        RECT 48.400 32.300 48.900 32.800 ;
        RECT 48.400 30.300 48.600 32.300 ;
        RECT 57.800 31.800 58.000 33.700 ;
        RECT 57.500 31.300 58.000 31.800 ;
        RECT 48.400 29.800 48.900 30.300 ;
        RECT 48.400 27.900 48.600 29.800 ;
        RECT 57.800 29.300 58.000 31.300 ;
        RECT 58.200 34.600 58.700 35.100 ;
        RECT 58.200 30.200 58.400 34.600 ;
        RECT 68.100 33.100 68.300 38.500 ;
        RECT 67.800 32.600 68.300 33.100 ;
        RECT 68.100 30.700 68.300 32.600 ;
        RECT 67.800 30.200 68.300 30.700 ;
        RECT 58.200 29.700 58.700 30.200 ;
        RECT 57.500 28.800 58.000 29.300 ;
        RECT 48.400 27.400 48.900 27.900 ;
        RECT 48.400 25.400 48.600 27.400 ;
        RECT 57.800 26.900 58.000 28.800 ;
        RECT 57.500 26.400 58.000 26.900 ;
        RECT 7.220 24.800 7.720 25.100 ;
        RECT 9.720 24.800 10.220 25.100 ;
        RECT 15.620 24.800 16.120 25.100 ;
        RECT 18.020 24.800 18.520 25.100 ;
        RECT 24.020 24.400 24.520 25.100 ;
        RECT 26.420 24.400 26.920 25.100 ;
        RECT 28.820 24.400 29.320 25.100 ;
        RECT 31.220 24.400 31.720 25.100 ;
        RECT 33.420 24.800 33.920 25.100 ;
        RECT 48.400 24.900 48.900 25.400 ;
        RECT 48.400 23.000 48.600 24.900 ;
        RECT 57.800 24.500 58.000 26.400 ;
        RECT 68.100 24.700 68.300 30.200 ;
        RECT 68.500 36.100 69.000 36.600 ;
        RECT 68.500 27.900 68.700 36.100 ;
        RECT 68.500 27.400 69.000 27.900 ;
        RECT 57.500 24.000 58.000 24.500 ;
        RECT 67.400 24.200 68.300 24.700 ;
        RECT 38.020 22.800 42.920 23.000 ;
        RECT 38.020 22.500 38.520 22.800 ;
        RECT 42.720 18.000 42.920 22.800 ;
        RECT 48.400 22.500 48.900 23.000 ;
        RECT 48.400 20.700 48.600 22.500 ;
        RECT 57.800 22.100 58.000 24.000 ;
        RECT 68.100 22.300 68.300 24.200 ;
        RECT 57.500 21.600 58.000 22.100 ;
        RECT 67.400 21.800 68.300 22.300 ;
        RECT 48.400 20.200 48.900 20.700 ;
        RECT 42.420 17.500 42.920 18.000 ;
        RECT 42.420 16.600 42.920 17.100 ;
        RECT 13.620 15.400 14.120 15.700 ;
        RECT 18.520 15.400 19.020 15.700 ;
        RECT 13.620 15.200 19.020 15.400 ;
        RECT 42.720 15.000 42.920 16.600 ;
        RECT 7.220 14.800 42.920 15.000 ;
        RECT 7.220 14.500 7.720 14.800 ;
        RECT 9.620 14.500 10.120 14.800 ;
        RECT 12.020 14.500 12.520 14.800 ;
        RECT 14.520 14.500 15.020 14.800 ;
        RECT 16.920 14.500 17.420 14.800 ;
        RECT 19.420 14.500 19.920 14.800 ;
        RECT 21.820 14.500 22.320 14.800 ;
        RECT 24.220 14.500 24.720 14.800 ;
        RECT 26.620 14.500 27.120 14.800 ;
        RECT 42.520 13.000 43.020 13.500 ;
        RECT 42.820 12.200 43.020 13.000 ;
        RECT 38.120 12.000 43.020 12.200 ;
        RECT 38.120 11.700 38.620 12.000 ;
        RECT 37.420 10.700 37.920 11.200 ;
        RECT 37.720 8.900 37.920 10.700 ;
        RECT 38.420 10.000 38.620 11.700 ;
        RECT 49.000 11.000 49.500 11.300 ;
        RECT 51.400 11.000 51.900 11.300 ;
        RECT 53.700 11.000 54.200 11.300 ;
        RECT 49.000 10.800 54.200 11.000 ;
        RECT 50.200 10.300 50.700 10.600 ;
        RECT 52.500 10.300 53.000 10.600 ;
        RECT 54.700 10.300 55.200 10.600 ;
        RECT 50.200 10.100 55.200 10.300 ;
        RECT 38.120 9.500 38.620 10.000 ;
        RECT 37.420 8.400 37.920 8.900 ;
        RECT 37.720 6.500 37.920 8.400 ;
        RECT 38.420 7.700 38.620 9.500 ;
        RECT 38.120 7.200 38.620 7.700 ;
        RECT 37.420 6.000 37.920 6.500 ;
        RECT 5.300 5.900 6.000 6.000 ;
        RECT 55.000 5.900 55.200 10.100 ;
        RECT 56.000 5.900 56.500 6.200 ;
        RECT 5.300 5.600 6.720 5.900 ;
        RECT 8.720 5.600 9.220 5.900 ;
        RECT 11.120 5.600 11.620 5.900 ;
        RECT 13.520 5.600 14.020 5.900 ;
        RECT 15.920 5.600 16.420 5.900 ;
        RECT 18.420 5.600 18.920 5.900 ;
        RECT 20.820 5.600 21.320 5.900 ;
        RECT 23.320 5.600 23.820 5.900 ;
        RECT 25.720 5.600 26.220 5.900 ;
        RECT 28.020 5.600 28.520 5.900 ;
        RECT 55.000 5.700 56.500 5.900 ;
        RECT 57.800 6.000 58.000 21.600 ;
        RECT 68.100 19.900 68.300 21.800 ;
        RECT 67.400 19.400 68.300 19.900 ;
        RECT 68.100 17.500 68.300 19.400 ;
        RECT 67.400 17.000 68.300 17.500 ;
        RECT 68.100 15.300 68.300 17.000 ;
        RECT 67.800 14.800 68.300 15.300 ;
        RECT 68.500 16.300 69.000 16.800 ;
        RECT 68.500 15.300 68.700 16.300 ;
        RECT 68.500 14.800 69.000 15.300 ;
        RECT 65.500 10.200 66.000 10.700 ;
        RECT 59.600 6.000 60.100 6.300 ;
        RECT 57.800 5.800 60.100 6.000 ;
        RECT 60.500 6.000 61.000 6.300 ;
        RECT 65.800 6.000 66.000 10.200 ;
        RECT 68.100 7.200 68.800 7.900 ;
        RECT 68.100 6.200 68.800 6.900 ;
        RECT 60.500 5.800 66.000 6.000 ;
        RECT 5.300 5.400 28.520 5.600 ;
        RECT 5.300 5.300 6.000 5.400 ;
        RECT 71.000 5.000 73.000 42.700 ;
        RECT 74.400 42.700 99.000 42.900 ;
        RECT 74.400 42.500 74.600 42.700 ;
        RECT 74.400 42.000 74.900 42.500 ;
        RECT 74.400 40.000 74.600 42.000 ;
        RECT 83.500 41.000 84.000 41.500 ;
        RECT 93.800 41.000 94.300 41.500 ;
        RECT 74.400 39.500 74.900 40.000 ;
        RECT 74.400 37.600 74.600 39.500 ;
        RECT 83.800 39.100 84.000 41.000 ;
        RECT 83.500 38.600 84.000 39.100 ;
        RECT 94.100 39.000 94.300 41.000 ;
        RECT 74.400 37.100 74.900 37.600 ;
        RECT 74.400 35.200 74.600 37.100 ;
        RECT 83.800 36.700 84.000 38.600 ;
        RECT 93.800 38.500 94.300 39.000 ;
        RECT 83.500 36.200 84.000 36.700 ;
        RECT 74.400 34.700 74.900 35.200 ;
        RECT 74.400 32.800 74.600 34.700 ;
        RECT 83.800 34.200 84.000 36.200 ;
        RECT 83.500 33.700 84.000 34.200 ;
        RECT 74.400 32.300 74.900 32.800 ;
        RECT 74.400 30.300 74.600 32.300 ;
        RECT 83.800 31.800 84.000 33.700 ;
        RECT 83.500 31.300 84.000 31.800 ;
        RECT 74.400 29.800 74.900 30.300 ;
        RECT 74.400 27.900 74.600 29.800 ;
        RECT 83.800 29.300 84.000 31.300 ;
        RECT 84.200 34.600 84.700 35.100 ;
        RECT 84.200 30.200 84.400 34.600 ;
        RECT 94.100 33.100 94.300 38.500 ;
        RECT 93.800 32.600 94.300 33.100 ;
        RECT 94.100 30.700 94.300 32.600 ;
        RECT 93.800 30.200 94.300 30.700 ;
        RECT 84.200 29.700 84.700 30.200 ;
        RECT 83.500 28.800 84.000 29.300 ;
        RECT 74.400 27.400 74.900 27.900 ;
        RECT 74.400 25.400 74.600 27.400 ;
        RECT 83.800 26.900 84.000 28.800 ;
        RECT 83.500 26.400 84.000 26.900 ;
        RECT 74.400 24.900 74.900 25.400 ;
        RECT 74.400 23.000 74.600 24.900 ;
        RECT 83.800 24.500 84.000 26.400 ;
        RECT 94.100 24.700 94.300 30.200 ;
        RECT 94.500 36.100 95.000 36.600 ;
        RECT 94.500 27.900 94.700 36.100 ;
        RECT 94.500 27.400 95.000 27.900 ;
        RECT 83.500 24.000 84.000 24.500 ;
        RECT 93.400 24.200 94.300 24.700 ;
        RECT 74.400 22.500 74.900 23.000 ;
        RECT 74.400 20.700 74.600 22.500 ;
        RECT 83.800 22.100 84.000 24.000 ;
        RECT 94.100 22.300 94.300 24.200 ;
        RECT 83.500 21.600 84.000 22.100 ;
        RECT 93.400 21.800 94.300 22.300 ;
        RECT 74.400 20.200 74.900 20.700 ;
        RECT 75.000 11.000 75.500 11.300 ;
        RECT 77.400 11.000 77.900 11.300 ;
        RECT 79.700 11.000 80.200 11.300 ;
        RECT 75.000 10.800 80.200 11.000 ;
        RECT 76.200 10.300 76.700 10.600 ;
        RECT 78.500 10.300 79.000 10.600 ;
        RECT 80.700 10.300 81.200 10.600 ;
        RECT 76.200 10.100 81.200 10.300 ;
        RECT 81.000 5.900 81.200 10.100 ;
        RECT 82.000 5.900 82.500 6.200 ;
        RECT 81.000 5.700 82.500 5.900 ;
        RECT 83.800 6.000 84.000 21.600 ;
        RECT 94.100 19.900 94.300 21.800 ;
        RECT 93.400 19.400 94.300 19.900 ;
        RECT 94.100 17.500 94.300 19.400 ;
        RECT 93.400 17.000 94.300 17.500 ;
        RECT 94.100 15.300 94.300 17.000 ;
        RECT 93.800 14.800 94.300 15.300 ;
        RECT 94.500 16.300 95.000 16.800 ;
        RECT 94.500 15.300 94.700 16.300 ;
        RECT 94.500 14.800 95.000 15.300 ;
        RECT 91.500 10.200 92.000 10.700 ;
        RECT 85.600 6.000 86.100 6.300 ;
        RECT 83.800 5.800 86.100 6.000 ;
        RECT 86.500 6.000 87.000 6.300 ;
        RECT 91.800 6.000 92.000 10.200 ;
        RECT 94.100 7.200 94.800 7.900 ;
        RECT 94.100 6.200 94.800 6.900 ;
        RECT 86.500 5.800 92.000 6.000 ;
        RECT 97.000 5.000 99.000 42.700 ;
        RECT 151.800 1.300 152.500 2.000 ;
      LAYER met3 ;
        RECT 96.800 223.700 97.500 224.400 ;
        RECT 99.600 223.700 100.300 224.400 ;
        RECT 102.300 223.700 103.000 224.400 ;
        RECT 105.100 223.700 105.800 224.400 ;
        RECT 107.900 223.700 108.600 224.400 ;
        RECT 110.700 223.700 111.400 224.400 ;
        RECT 113.400 223.700 114.100 224.400 ;
        RECT 116.100 223.700 116.800 224.400 ;
        RECT 118.900 223.700 119.600 224.400 ;
        RECT 121.700 223.700 122.400 224.400 ;
        RECT 124.500 223.700 125.200 224.400 ;
        RECT 127.200 223.700 127.900 224.400 ;
        RECT 130.000 223.700 130.700 224.400 ;
        RECT 132.800 223.700 133.500 224.400 ;
        RECT 135.500 223.700 136.200 224.400 ;
        RECT 138.300 223.700 139.000 224.400 ;
        RECT 96.800 221.000 97.100 223.700 ;
        RECT 99.600 221.000 99.900 223.700 ;
        RECT 102.300 221.000 102.600 223.700 ;
        RECT 105.100 221.000 105.400 223.700 ;
        RECT 96.800 220.300 97.500 221.000 ;
        RECT 99.600 220.300 100.300 221.000 ;
        RECT 102.300 220.300 103.000 221.000 ;
        RECT 105.100 220.300 105.800 221.000 ;
        RECT 119.000 216.700 119.300 223.700 ;
        RECT 44.800 216.400 119.300 216.700 ;
        RECT 44.800 209.600 45.100 216.400 ;
        RECT 121.800 216.100 122.100 223.700 ;
        RECT 45.800 215.800 122.100 216.100 ;
        RECT 45.800 209.600 46.100 215.800 ;
        RECT 124.500 215.500 124.800 223.700 ;
        RECT 46.800 215.200 124.800 215.500 ;
        RECT 46.800 209.600 47.100 215.200 ;
        RECT 127.300 214.900 127.600 223.700 ;
        RECT 47.800 214.600 127.600 214.900 ;
        RECT 47.800 209.600 48.100 214.600 ;
        RECT 130.100 214.300 130.400 223.700 ;
        RECT 48.800 214.000 130.400 214.300 ;
        RECT 48.800 209.600 49.100 214.000 ;
        RECT 132.900 213.700 133.200 223.700 ;
        RECT 49.800 213.400 133.200 213.700 ;
        RECT 49.800 209.600 50.100 213.400 ;
        RECT 135.600 213.100 135.900 223.700 ;
        RECT 50.800 212.800 135.900 213.100 ;
        RECT 50.800 209.600 51.300 212.800 ;
        RECT 138.300 212.500 138.600 223.700 ;
        RECT 51.800 212.200 138.600 212.500 ;
        RECT 51.800 209.600 52.100 212.200 ;
        RECT 44.800 209.400 45.400 209.600 ;
        RECT 45.800 209.400 46.400 209.600 ;
        RECT 46.800 209.400 47.400 209.600 ;
        RECT 47.800 209.400 48.400 209.600 ;
        RECT 48.800 209.400 49.400 209.600 ;
        RECT 49.800 209.400 50.400 209.600 ;
        RECT 50.800 209.400 51.400 209.600 ;
        RECT 51.800 209.400 52.400 209.600 ;
        RECT 44.900 209.100 45.400 209.400 ;
        RECT 45.900 209.100 46.400 209.400 ;
        RECT 46.900 209.100 47.400 209.400 ;
        RECT 47.900 209.100 48.400 209.400 ;
        RECT 48.900 209.100 49.400 209.400 ;
        RECT 49.900 209.100 50.400 209.400 ;
        RECT 50.900 209.100 51.400 209.400 ;
        RECT 51.900 209.100 52.400 209.400 ;
        RECT 2.300 207.700 3.000 208.400 ;
        RECT 40.900 207.100 41.600 207.800 ;
        RECT 41.900 207.100 42.600 207.800 ;
        RECT 5.300 187.300 6.000 188.000 ;
        RECT 2.300 181.700 3.000 182.400 ;
        RECT 40.900 181.100 41.600 181.800 ;
        RECT 41.900 181.100 42.600 181.800 ;
        RECT 5.300 161.300 6.000 162.000 ;
        RECT 2.300 155.700 3.000 156.400 ;
        RECT 40.900 155.100 41.600 155.800 ;
        RECT 41.900 155.100 42.600 155.800 ;
        RECT 5.300 135.300 6.000 136.000 ;
        RECT 68.100 133.200 68.800 133.900 ;
        RECT 94.100 133.200 94.800 133.900 ;
        RECT 68.100 132.200 68.800 132.900 ;
        RECT 94.100 132.200 94.800 132.900 ;
        RECT 2.300 129.700 3.000 130.400 ;
        RECT 40.900 129.100 41.600 129.800 ;
        RECT 41.900 129.100 42.600 129.800 ;
        RECT 5.300 109.300 6.000 110.000 ;
        RECT 2.300 103.700 3.000 104.400 ;
        RECT 40.900 103.100 41.600 103.800 ;
        RECT 41.900 103.100 42.600 103.800 ;
        RECT 68.100 91.200 68.800 91.900 ;
        RECT 94.100 91.200 94.800 91.900 ;
        RECT 68.100 90.200 68.800 90.900 ;
        RECT 94.100 90.200 94.800 90.900 ;
        RECT 5.300 83.300 6.000 84.000 ;
        RECT 2.300 77.700 3.000 78.400 ;
        RECT 40.900 77.100 41.600 77.800 ;
        RECT 41.900 77.100 42.600 77.800 ;
        RECT 5.300 57.300 6.000 58.000 ;
        RECT 2.300 51.700 3.000 52.400 ;
        RECT 40.900 51.100 41.600 51.800 ;
        RECT 41.900 51.100 42.600 51.800 ;
        RECT 68.100 49.200 68.800 49.900 ;
        RECT 94.100 49.200 94.800 49.900 ;
        RECT 68.100 48.200 68.800 48.900 ;
        RECT 94.100 48.200 94.800 48.900 ;
        RECT 5.300 31.300 6.000 32.000 ;
        RECT 2.300 25.700 3.000 26.400 ;
        RECT 40.900 25.100 41.600 25.800 ;
        RECT 41.900 25.100 42.600 25.800 ;
        RECT 68.100 7.200 68.800 7.900 ;
        RECT 94.100 7.200 94.800 7.900 ;
        RECT 68.100 6.200 68.800 6.900 ;
        RECT 94.100 6.200 94.800 6.900 ;
        RECT 5.300 5.300 6.000 6.000 ;
        RECT 151.800 1.300 152.500 2.000 ;
      LAYER met4 ;
        RECT 30.970 224.760 31.000 225.100 ;
        RECT 33.730 224.760 33.800 225.100 ;
        RECT 36.490 224.760 36.500 225.100 ;
        RECT 39.250 224.760 39.300 225.100 ;
        RECT 30.700 224.400 31.000 224.760 ;
        RECT 33.500 224.400 33.800 224.760 ;
        RECT 36.200 224.400 36.500 224.760 ;
        RECT 39.000 224.400 39.300 224.760 ;
        RECT 41.700 224.760 41.710 225.100 ;
        RECT 44.770 224.760 44.800 225.100 ;
        RECT 47.530 224.760 47.600 225.100 ;
        RECT 50.290 224.760 50.300 225.100 ;
        RECT 53.050 224.760 53.100 225.100 ;
        RECT 41.700 224.400 42.000 224.760 ;
        RECT 44.500 224.400 44.800 224.760 ;
        RECT 47.300 224.400 47.600 224.760 ;
        RECT 50.000 224.400 50.300 224.760 ;
        RECT 52.800 224.400 53.100 224.760 ;
        RECT 55.500 224.760 55.510 225.100 ;
        RECT 58.570 224.760 58.600 225.100 ;
        RECT 61.330 224.760 61.400 225.100 ;
        RECT 64.090 224.760 64.100 225.100 ;
        RECT 66.850 224.760 66.900 225.100 ;
        RECT 55.500 224.400 55.800 224.760 ;
        RECT 58.300 224.400 58.600 224.760 ;
        RECT 61.100 224.400 61.400 224.760 ;
        RECT 63.800 224.400 64.100 224.760 ;
        RECT 66.600 224.400 66.900 224.760 ;
        RECT 69.300 224.760 69.310 225.100 ;
        RECT 72.370 224.760 72.400 225.100 ;
        RECT 75.130 224.760 75.200 225.100 ;
        RECT 77.890 224.760 77.900 225.100 ;
        RECT 80.650 224.760 80.700 225.100 ;
        RECT 69.300 224.400 69.600 224.760 ;
        RECT 72.100 224.400 72.400 224.760 ;
        RECT 74.900 224.400 75.200 224.760 ;
        RECT 77.600 224.400 77.900 224.760 ;
        RECT 80.400 224.400 80.700 224.760 ;
        RECT 83.100 224.760 83.110 225.100 ;
        RECT 86.170 224.760 86.200 225.100 ;
        RECT 83.100 224.400 83.400 224.760 ;
        RECT 85.900 224.400 86.200 224.760 ;
        RECT 88.600 224.760 88.630 225.100 ;
        RECT 91.690 224.760 91.700 225.100 ;
        RECT 94.450 224.760 94.500 225.100 ;
        RECT 88.600 224.400 88.900 224.760 ;
        RECT 91.400 224.400 91.700 224.760 ;
        RECT 94.200 224.400 94.500 224.760 ;
        RECT 96.900 224.760 96.910 224.900 ;
        RECT 99.970 224.760 100.000 224.900 ;
        RECT 96.900 224.400 97.200 224.760 ;
        RECT 99.700 224.400 100.000 224.760 ;
        RECT 102.400 224.760 102.430 224.900 ;
        RECT 105.490 224.760 105.500 224.900 ;
        RECT 102.400 224.400 102.700 224.760 ;
        RECT 105.200 224.400 105.500 224.760 ;
        RECT 107.900 224.760 107.950 224.900 ;
        RECT 108.250 224.760 108.300 224.900 ;
        RECT 107.900 224.400 108.300 224.760 ;
        RECT 110.700 224.760 110.710 224.900 ;
        RECT 113.770 224.760 113.800 225.000 ;
        RECT 110.700 224.400 111.000 224.760 ;
        RECT 113.500 224.400 113.800 224.760 ;
        RECT 116.200 224.760 116.230 225.000 ;
        RECT 118.900 224.760 118.990 225.000 ;
        RECT 121.700 224.760 121.750 225.000 ;
        RECT 124.500 224.760 124.510 225.000 ;
        RECT 127.200 224.760 127.270 225.000 ;
        RECT 130.000 224.760 130.030 225.000 ;
        RECT 133.090 224.760 133.100 225.000 ;
        RECT 116.200 224.400 116.500 224.760 ;
        RECT 118.900 224.400 119.200 224.760 ;
        RECT 121.700 224.400 122.000 224.760 ;
        RECT 124.500 224.400 124.800 224.760 ;
        RECT 127.200 224.400 127.500 224.760 ;
        RECT 130.000 224.400 130.300 224.760 ;
        RECT 132.800 224.400 133.100 224.760 ;
        RECT 135.500 224.760 135.550 225.000 ;
        RECT 138.300 224.760 138.310 225.000 ;
        RECT 135.500 224.400 135.800 224.760 ;
        RECT 138.300 224.400 138.600 224.760 ;
        RECT 6.300 224.100 94.500 224.400 ;
        RECT 6.300 220.800 6.600 224.100 ;
        RECT 96.800 223.700 97.500 224.400 ;
        RECT 99.600 223.700 100.300 224.400 ;
        RECT 102.300 223.700 103.000 224.400 ;
        RECT 105.100 223.700 105.800 224.400 ;
        RECT 107.900 223.700 108.600 224.400 ;
        RECT 110.700 223.700 111.400 224.400 ;
        RECT 113.400 223.700 114.100 224.400 ;
        RECT 116.100 223.700 116.800 224.400 ;
        RECT 118.900 223.700 119.600 224.400 ;
        RECT 121.700 223.700 122.400 224.400 ;
        RECT 124.500 223.700 125.200 224.400 ;
        RECT 127.200 223.700 127.900 224.400 ;
        RECT 130.000 223.700 130.700 224.400 ;
        RECT 132.800 223.700 133.500 224.400 ;
        RECT 135.500 223.700 136.200 224.400 ;
        RECT 138.300 223.700 139.000 224.400 ;
        RECT 107.900 223.400 108.200 223.700 ;
        RECT 5.700 220.760 6.600 220.800 ;
        RECT 6.000 220.500 6.600 220.760 ;
        RECT 70.900 223.100 108.200 223.400 ;
        RECT 40.900 207.400 41.600 207.800 ;
        RECT 41.900 207.400 42.600 207.800 ;
        RECT 40.900 207.100 42.600 207.400 ;
        RECT 40.900 181.400 41.600 181.800 ;
        RECT 41.900 181.400 42.600 181.800 ;
        RECT 40.900 181.100 42.600 181.400 ;
        RECT 40.900 155.400 41.600 155.800 ;
        RECT 41.900 155.400 42.600 155.800 ;
        RECT 40.900 155.100 42.600 155.400 ;
        RECT 68.100 133.200 68.800 133.900 ;
        RECT 68.100 132.900 68.400 133.200 ;
        RECT 68.100 132.500 68.800 132.900 ;
        RECT 70.900 132.500 71.200 223.100 ;
        RECT 110.700 222.800 111.000 223.700 ;
        RECT 68.100 132.200 71.200 132.500 ;
        RECT 71.500 222.500 111.000 222.800 ;
        RECT 40.900 129.400 41.600 129.800 ;
        RECT 41.900 129.400 42.600 129.800 ;
        RECT 40.900 129.100 42.600 129.400 ;
        RECT 40.900 103.400 41.600 103.800 ;
        RECT 41.900 103.400 42.600 103.800 ;
        RECT 40.900 103.100 42.600 103.400 ;
        RECT 68.100 91.200 68.800 91.900 ;
        RECT 68.100 90.900 68.400 91.200 ;
        RECT 68.100 90.500 68.800 90.900 ;
        RECT 71.500 90.500 71.800 222.500 ;
        RECT 113.400 222.200 113.700 223.700 ;
        RECT 68.100 90.200 71.800 90.500 ;
        RECT 72.100 221.900 113.700 222.200 ;
        RECT 40.900 77.400 41.600 77.800 ;
        RECT 41.900 77.400 42.600 77.800 ;
        RECT 40.900 77.100 42.600 77.400 ;
        RECT 40.900 51.400 41.600 51.800 ;
        RECT 41.900 51.400 42.600 51.800 ;
        RECT 40.900 51.100 42.600 51.400 ;
        RECT 68.100 49.200 68.800 49.900 ;
        RECT 68.100 48.900 68.400 49.200 ;
        RECT 68.100 48.500 68.800 48.900 ;
        RECT 72.100 48.500 72.400 221.900 ;
        RECT 116.100 221.600 116.400 223.700 ;
        RECT 68.100 48.200 72.400 48.500 ;
        RECT 72.700 221.300 116.400 221.600 ;
        RECT 40.900 25.400 41.600 25.800 ;
        RECT 41.900 25.400 42.600 25.800 ;
        RECT 40.900 25.100 42.600 25.400 ;
        RECT 68.100 7.200 68.800 7.900 ;
        RECT 68.100 6.900 68.400 7.200 ;
        RECT 68.100 6.500 68.800 6.900 ;
        RECT 72.700 6.500 73.000 221.300 ;
        RECT 96.800 220.300 97.500 221.000 ;
        RECT 99.600 220.300 100.300 221.000 ;
        RECT 102.300 220.300 103.000 221.000 ;
        RECT 105.100 220.300 105.800 221.000 ;
        RECT 94.100 133.200 94.800 133.900 ;
        RECT 94.100 132.900 94.400 133.200 ;
        RECT 94.100 132.500 94.800 132.900 ;
        RECT 96.900 132.500 97.200 220.300 ;
        RECT 99.600 220.000 99.900 220.300 ;
        RECT 94.100 132.200 97.200 132.500 ;
        RECT 97.500 219.700 99.900 220.000 ;
        RECT 94.100 91.200 94.800 91.900 ;
        RECT 94.100 90.900 94.400 91.200 ;
        RECT 94.100 90.500 94.800 90.900 ;
        RECT 97.500 90.500 97.800 219.700 ;
        RECT 102.300 219.400 102.600 220.300 ;
        RECT 94.100 90.200 97.800 90.500 ;
        RECT 98.100 219.100 102.600 219.400 ;
        RECT 94.100 49.200 94.800 49.900 ;
        RECT 94.100 48.900 94.400 49.200 ;
        RECT 94.100 48.500 94.800 48.900 ;
        RECT 98.100 48.500 98.400 219.100 ;
        RECT 105.100 218.800 105.400 220.300 ;
        RECT 94.100 48.200 98.400 48.500 ;
        RECT 98.700 218.500 105.400 218.800 ;
        RECT 68.100 6.200 73.000 6.500 ;
        RECT 94.100 7.200 94.800 7.900 ;
        RECT 94.100 6.900 94.400 7.200 ;
        RECT 94.100 6.500 94.800 6.900 ;
        RECT 98.700 6.500 99.000 218.500 ;
        RECT 94.100 6.200 99.000 6.500 ;
        RECT 151.800 1.300 152.500 2.000 ;
        RECT 151.800 1.000 152.100 1.300 ;
        RECT 151.800 0.700 151.810 1.000 ;
  END
END tt_um_rburt16_bias_generator
END LIBRARY

