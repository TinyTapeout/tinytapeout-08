module test_tt;
  initial begin
    $display("Hello from test_tt!");
    $finish;
  end
endmodule
