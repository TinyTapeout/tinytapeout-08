VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_a1k0n_demo
  CLASS BLOCK ;
  FOREIGN tt_um_a1k0n_demo ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.450 2.480 62.050 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.320 2.480 100.920 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.190 2.480 139.790 223.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.150 2.480 58.750 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.020 2.480 97.620 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.890 2.480 136.490 223.280 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 158.240 223.125 ;
      LAYER met1 ;
        RECT 0.070 0.040 160.930 225.720 ;
      LAYER met2 ;
        RECT 0.090 0.010 160.900 225.750 ;
      LAYER met3 ;
        RECT 0.065 1.535 160.475 225.585 ;
      LAYER met4 ;
        RECT 3.975 224.360 30.270 224.905 ;
        RECT 31.370 224.360 33.030 224.905 ;
        RECT 34.130 224.360 35.790 224.905 ;
        RECT 36.890 224.360 38.550 224.905 ;
        RECT 39.650 224.360 41.310 224.905 ;
        RECT 42.410 224.360 44.070 224.905 ;
        RECT 45.170 224.360 46.830 224.905 ;
        RECT 47.930 224.360 49.590 224.905 ;
        RECT 50.690 224.360 52.350 224.905 ;
        RECT 53.450 224.360 55.110 224.905 ;
        RECT 56.210 224.360 57.870 224.905 ;
        RECT 58.970 224.360 60.630 224.905 ;
        RECT 61.730 224.360 63.390 224.905 ;
        RECT 64.490 224.360 66.150 224.905 ;
        RECT 67.250 224.360 68.910 224.905 ;
        RECT 70.010 224.360 71.670 224.905 ;
        RECT 72.770 224.360 74.430 224.905 ;
        RECT 75.530 224.360 77.190 224.905 ;
        RECT 78.290 224.360 79.950 224.905 ;
        RECT 81.050 224.360 82.710 224.905 ;
        RECT 83.810 224.360 85.470 224.905 ;
        RECT 86.570 224.360 88.230 224.905 ;
        RECT 89.330 224.360 90.990 224.905 ;
        RECT 92.090 224.360 93.750 224.905 ;
        RECT 94.850 224.360 96.510 224.905 ;
        RECT 97.610 224.360 99.270 224.905 ;
        RECT 100.370 224.360 102.030 224.905 ;
        RECT 103.130 224.360 104.790 224.905 ;
        RECT 105.890 224.360 107.550 224.905 ;
        RECT 108.650 224.360 110.310 224.905 ;
        RECT 111.410 224.360 113.070 224.905 ;
        RECT 114.170 224.360 115.830 224.905 ;
        RECT 116.930 224.360 118.590 224.905 ;
        RECT 119.690 224.360 121.350 224.905 ;
        RECT 122.450 224.360 124.110 224.905 ;
        RECT 125.210 224.360 126.870 224.905 ;
        RECT 127.970 224.360 129.630 224.905 ;
        RECT 130.730 224.360 132.390 224.905 ;
        RECT 133.490 224.360 135.150 224.905 ;
        RECT 136.250 224.360 137.910 224.905 ;
        RECT 139.010 224.360 140.670 224.905 ;
        RECT 141.770 224.360 143.430 224.905 ;
        RECT 144.530 224.360 146.190 224.905 ;
        RECT 147.290 224.360 151.505 224.905 ;
        RECT 3.975 223.680 151.505 224.360 ;
        RECT 3.975 2.080 17.880 223.680 ;
        RECT 20.280 2.080 21.180 223.680 ;
        RECT 23.580 2.080 56.750 223.680 ;
        RECT 59.150 2.080 60.050 223.680 ;
        RECT 62.450 2.080 95.620 223.680 ;
        RECT 98.020 2.080 98.920 223.680 ;
        RECT 101.320 2.080 134.490 223.680 ;
        RECT 136.890 2.080 137.790 223.680 ;
        RECT 140.190 2.080 151.505 223.680 ;
        RECT 3.975 1.535 151.505 2.080 ;
  END
END tt_um_a1k0n_demo
END LIBRARY

