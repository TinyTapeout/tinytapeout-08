module tt_um_ran_DanielZhu (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input VPWR;
 input VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire clknet_0_clk;
 wire \tt_16bitran.connection[0] ;
 wire \tt_16bitran.connection[10] ;
 wire \tt_16bitran.connection[11] ;
 wire \tt_16bitran.connection[12] ;
 wire \tt_16bitran.connection[13] ;
 wire \tt_16bitran.connection[14] ;
 wire \tt_16bitran.connection[15] ;
 wire \tt_16bitran.connection[16] ;
 wire \tt_16bitran.connection[1] ;
 wire \tt_16bitran.connection[2] ;
 wire \tt_16bitran.connection[3] ;
 wire \tt_16bitran.connection[4] ;
 wire \tt_16bitran.connection[5] ;
 wire \tt_16bitran.connection[6] ;
 wire \tt_16bitran.connection[7] ;
 wire \tt_16bitran.connection[8] ;
 wire \tt_16bitran.connection[9] ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.key ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.key ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.key ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.key ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[0].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[0].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[1].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[1].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[2].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[2].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[3].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[3].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[4].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[4].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[5].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[5].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[6].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[6].multblock.nand_gate_2.B_1 ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.a ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.b ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.c ;
 wire \tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.d ;
 wire \tt_finalprocess.genblk1[7].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[7].multblock.nand_gate_2.B_1 ;
 wire \tt_invring1.ringosc1[0].inv.a ;
 wire \tt_invring1.ringosc1[0].inv.y ;
 wire \tt_invring1.ringosc1[10].inv.a ;
 wire \tt_invring1.ringosc1[10].inv.y ;
 wire \tt_invring1.ringosc1[1].inv.y ;
 wire \tt_invring1.ringosc1[2].inv.y ;
 wire \tt_invring1.ringosc1[3].inv.y ;
 wire \tt_invring1.ringosc1[4].inv.y ;
 wire \tt_invring1.ringosc1[5].inv.y ;
 wire \tt_invring1.ringosc1[6].inv.y ;
 wire \tt_invring1.ringosc1[7].inv.y ;
 wire \tt_invring1.ringosc1[8].inv.y ;
 wire \tt_invring1.ringosc2[0].inv.a ;
 wire \tt_invring1.ringosc2[0].inv.y ;
 wire \tt_invring1.ringosc2[10].inv.a ;
 wire \tt_invring1.ringosc2[10].inv.y ;
 wire \tt_invring1.ringosc2[11].inv.y ;
 wire \tt_invring1.ringosc2[12].inv.y ;
 wire \tt_invring1.ringosc2[13].inv.y ;
 wire \tt_invring1.ringosc2[14].inv.y ;
 wire \tt_invring1.ringosc2[15].inv.y ;
 wire \tt_invring1.ringosc2[16].inv.y ;
 wire \tt_invring1.ringosc2[17].inv.y ;
 wire \tt_invring1.ringosc2[18].inv.y ;
 wire \tt_invring1.ringosc2[1].inv.y ;
 wire \tt_invring1.ringosc2[2].inv.y ;
 wire \tt_invring1.ringosc2[3].inv.y ;
 wire \tt_invring1.ringosc2[4].inv.y ;
 wire \tt_invring1.ringosc2[5].inv.y ;
 wire \tt_invring1.ringosc2[6].inv.y ;
 wire \tt_invring1.ringosc2[7].inv.y ;
 wire \tt_invring1.ringosc2[8].inv.y ;
 wire \tt_invring1.ringosc3[0].inv.a ;
 wire \tt_invring1.ringosc3[0].inv.y ;
 wire \tt_invring1.ringosc3[10].inv.a ;
 wire \tt_invring1.ringosc3[10].inv.y ;
 wire \tt_invring1.ringosc3[11].inv.y ;
 wire \tt_invring1.ringosc3[12].inv.y ;
 wire \tt_invring1.ringosc3[13].inv.y ;
 wire \tt_invring1.ringosc3[14].inv.y ;
 wire \tt_invring1.ringosc3[15].inv.y ;
 wire \tt_invring1.ringosc3[16].inv.y ;
 wire \tt_invring1.ringosc3[17].inv.y ;
 wire \tt_invring1.ringosc3[18].inv.y ;
 wire \tt_invring1.ringosc3[19].inv.y ;
 wire \tt_invring1.ringosc3[1].inv.y ;
 wire \tt_invring1.ringosc3[20].inv.y ;
 wire \tt_invring1.ringosc3[21].inv.y ;
 wire \tt_invring1.ringosc3[22].inv.y ;
 wire \tt_invring1.ringosc3[2].inv.y ;
 wire \tt_invring1.ringosc3[3].inv.y ;
 wire \tt_invring1.ringosc3[4].inv.y ;
 wire \tt_invring1.ringosc3[5].inv.y ;
 wire \tt_invring1.ringosc3[6].inv.y ;
 wire \tt_invring1.ringosc3[7].inv.y ;
 wire \tt_invring1.ringosc3[8].inv.y ;
 wire \tt_invring1.ringosc4[0].inv.a ;
 wire \tt_invring1.ringosc4[0].inv.y ;
 wire \tt_invring1.ringosc4[10].inv.a ;
 wire \tt_invring1.ringosc4[10].inv.y ;
 wire \tt_invring1.ringosc4[11].inv.y ;
 wire \tt_invring1.ringosc4[12].inv.y ;
 wire \tt_invring1.ringosc4[13].inv.y ;
 wire \tt_invring1.ringosc4[14].inv.y ;
 wire \tt_invring1.ringosc4[15].inv.y ;
 wire \tt_invring1.ringosc4[16].inv.y ;
 wire \tt_invring1.ringosc4[17].inv.y ;
 wire \tt_invring1.ringosc4[18].inv.y ;
 wire \tt_invring1.ringosc4[19].inv.y ;
 wire \tt_invring1.ringosc4[1].inv.y ;
 wire \tt_invring1.ringosc4[20].inv.y ;
 wire \tt_invring1.ringosc4[21].inv.y ;
 wire \tt_invring1.ringosc4[22].inv.y ;
 wire \tt_invring1.ringosc4[23].inv.y ;
 wire \tt_invring1.ringosc4[24].inv.y ;
 wire \tt_invring1.ringosc4[25].inv.y ;
 wire \tt_invring1.ringosc4[26].inv.y ;
 wire \tt_invring1.ringosc4[27].inv.y ;
 wire \tt_invring1.ringosc4[28].inv.y ;
 wire \tt_invring1.ringosc4[2].inv.y ;
 wire \tt_invring1.ringosc4[3].inv.y ;
 wire \tt_invring1.ringosc4[4].inv.y ;
 wire \tt_invring1.ringosc4[5].inv.y ;
 wire \tt_invring1.ringosc4[6].inv.y ;
 wire \tt_invring1.ringosc4[7].inv.y ;
 wire \tt_invring1.ringosc4[8].inv.y ;
 wire \tt_invring1.ringosc5[0].inv.a ;
 wire \tt_invring1.ringosc5[0].inv.y ;
 wire \tt_invring1.ringosc5[10].inv.a ;
 wire \tt_invring1.ringosc5[10].inv.y ;
 wire \tt_invring1.ringosc5[11].inv.y ;
 wire \tt_invring1.ringosc5[12].inv.y ;
 wire \tt_invring1.ringosc5[13].inv.y ;
 wire \tt_invring1.ringosc5[14].inv.y ;
 wire \tt_invring1.ringosc5[15].inv.y ;
 wire \tt_invring1.ringosc5[16].inv.y ;
 wire \tt_invring1.ringosc5[17].inv.y ;
 wire \tt_invring1.ringosc5[18].inv.y ;
 wire \tt_invring1.ringosc5[19].inv.y ;
 wire \tt_invring1.ringosc5[1].inv.y ;
 wire \tt_invring1.ringosc5[20].inv.y ;
 wire \tt_invring1.ringosc5[21].inv.y ;
 wire \tt_invring1.ringosc5[22].inv.y ;
 wire \tt_invring1.ringosc5[23].inv.y ;
 wire \tt_invring1.ringosc5[24].inv.y ;
 wire \tt_invring1.ringosc5[25].inv.y ;
 wire \tt_invring1.ringosc5[26].inv.y ;
 wire \tt_invring1.ringosc5[27].inv.y ;
 wire \tt_invring1.ringosc5[28].inv.y ;
 wire \tt_invring1.ringosc5[29].inv.y ;
 wire \tt_invring1.ringosc5[2].inv.y ;
 wire \tt_invring1.ringosc5[30].inv.y ;
 wire \tt_invring1.ringosc5[31].inv.y ;
 wire \tt_invring1.ringosc5[32].inv.y ;
 wire \tt_invring1.ringosc5[33].inv.y ;
 wire \tt_invring1.ringosc5[34].inv.y ;
 wire \tt_invring1.ringosc5[35].inv.y ;
 wire \tt_invring1.ringosc5[36].inv.y ;
 wire \tt_invring1.ringosc5[3].inv.y ;
 wire \tt_invring1.ringosc5[4].inv.y ;
 wire \tt_invring1.ringosc5[5].inv.y ;
 wire \tt_invring1.ringosc5[6].inv.y ;
 wire \tt_invring1.ringosc5[7].inv.y ;
 wire \tt_invring1.ringosc5[8].inv.y ;
 wire \tt_invring1.ringosc6[0].inv.a ;
 wire \tt_invring1.ringosc6[0].inv.y ;
 wire \tt_invring1.ringosc6[10].inv.a ;
 wire \tt_invring1.ringosc6[10].inv.y ;
 wire \tt_invring1.ringosc6[11].inv.y ;
 wire \tt_invring1.ringosc6[12].inv.y ;
 wire \tt_invring1.ringosc6[13].inv.y ;
 wire \tt_invring1.ringosc6[14].inv.y ;
 wire \tt_invring1.ringosc6[15].inv.y ;
 wire \tt_invring1.ringosc6[16].inv.y ;
 wire \tt_invring1.ringosc6[17].inv.y ;
 wire \tt_invring1.ringosc6[18].inv.y ;
 wire \tt_invring1.ringosc6[19].inv.y ;
 wire \tt_invring1.ringosc6[1].inv.y ;
 wire \tt_invring1.ringosc6[20].inv.y ;
 wire \tt_invring1.ringosc6[21].inv.y ;
 wire \tt_invring1.ringosc6[22].inv.y ;
 wire \tt_invring1.ringosc6[23].inv.y ;
 wire \tt_invring1.ringosc6[24].inv.y ;
 wire \tt_invring1.ringosc6[25].inv.y ;
 wire \tt_invring1.ringosc6[26].inv.y ;
 wire \tt_invring1.ringosc6[27].inv.y ;
 wire \tt_invring1.ringosc6[28].inv.y ;
 wire \tt_invring1.ringosc6[29].inv.y ;
 wire \tt_invring1.ringosc6[2].inv.y ;
 wire \tt_invring1.ringosc6[30].inv.y ;
 wire \tt_invring1.ringosc6[31].inv.y ;
 wire \tt_invring1.ringosc6[32].inv.y ;
 wire \tt_invring1.ringosc6[33].inv.y ;
 wire \tt_invring1.ringosc6[34].inv.y ;
 wire \tt_invring1.ringosc6[35].inv.y ;
 wire \tt_invring1.ringosc6[36].inv.y ;
 wire \tt_invring1.ringosc6[37].inv.y ;
 wire \tt_invring1.ringosc6[38].inv.y ;
 wire \tt_invring1.ringosc6[39].inv.y ;
 wire \tt_invring1.ringosc6[3].inv.y ;
 wire \tt_invring1.ringosc6[40].inv.y ;
 wire \tt_invring1.ringosc6[4].inv.y ;
 wire \tt_invring1.ringosc6[5].inv.y ;
 wire \tt_invring1.ringosc6[6].inv.y ;
 wire \tt_invring1.ringosc6[7].inv.y ;
 wire \tt_invring1.ringosc6[8].inv.y ;
 wire \tt_invring1.ringosc7[0].inv.a ;
 wire \tt_invring1.ringosc7[0].inv.y ;
 wire \tt_invring1.ringosc7[10].inv.a ;
 wire \tt_invring1.ringosc7[10].inv.y ;
 wire \tt_invring1.ringosc7[11].inv.y ;
 wire \tt_invring1.ringosc7[12].inv.y ;
 wire \tt_invring1.ringosc7[13].inv.y ;
 wire \tt_invring1.ringosc7[14].inv.y ;
 wire \tt_invring1.ringosc7[15].inv.y ;
 wire \tt_invring1.ringosc7[16].inv.y ;
 wire \tt_invring1.ringosc7[17].inv.y ;
 wire \tt_invring1.ringosc7[18].inv.y ;
 wire \tt_invring1.ringosc7[19].inv.y ;
 wire \tt_invring1.ringosc7[1].inv.y ;
 wire \tt_invring1.ringosc7[20].inv.y ;
 wire \tt_invring1.ringosc7[21].inv.y ;
 wire \tt_invring1.ringosc7[22].inv.y ;
 wire \tt_invring1.ringosc7[23].inv.y ;
 wire \tt_invring1.ringosc7[24].inv.y ;
 wire \tt_invring1.ringosc7[25].inv.y ;
 wire \tt_invring1.ringosc7[26].inv.y ;
 wire \tt_invring1.ringosc7[27].inv.y ;
 wire \tt_invring1.ringosc7[28].inv.y ;
 wire \tt_invring1.ringosc7[29].inv.y ;
 wire \tt_invring1.ringosc7[2].inv.y ;
 wire \tt_invring1.ringosc7[30].inv.y ;
 wire \tt_invring1.ringosc7[31].inv.y ;
 wire \tt_invring1.ringosc7[32].inv.y ;
 wire \tt_invring1.ringosc7[33].inv.y ;
 wire \tt_invring1.ringosc7[34].inv.y ;
 wire \tt_invring1.ringosc7[35].inv.y ;
 wire \tt_invring1.ringosc7[36].inv.y ;
 wire \tt_invring1.ringosc7[37].inv.y ;
 wire \tt_invring1.ringosc7[38].inv.y ;
 wire \tt_invring1.ringosc7[39].inv.y ;
 wire \tt_invring1.ringosc7[3].inv.y ;
 wire \tt_invring1.ringosc7[40].inv.y ;
 wire \tt_invring1.ringosc7[41].inv.y ;
 wire \tt_invring1.ringosc7[42].inv.y ;
 wire \tt_invring1.ringosc7[43].inv.y ;
 wire \tt_invring1.ringosc7[44].inv.y ;
 wire \tt_invring1.ringosc7[45].inv.y ;
 wire \tt_invring1.ringosc7[46].inv.y ;
 wire \tt_invring1.ringosc7[4].inv.y ;
 wire \tt_invring1.ringosc7[5].inv.y ;
 wire \tt_invring1.ringosc7[6].inv.y ;
 wire \tt_invring1.ringosc7[7].inv.y ;
 wire \tt_invring1.ringosc7[8].inv.y ;
 wire \tt_invring1.ringosc8[0].inv.a ;
 wire \tt_invring1.ringosc8[0].inv.y ;
 wire \tt_invring1.ringosc8[10].inv.a ;
 wire \tt_invring1.ringosc8[10].inv.y ;
 wire \tt_invring1.ringosc8[11].inv.y ;
 wire \tt_invring1.ringosc8[12].inv.y ;
 wire \tt_invring1.ringosc8[13].inv.y ;
 wire \tt_invring1.ringosc8[14].inv.y ;
 wire \tt_invring1.ringosc8[15].inv.y ;
 wire \tt_invring1.ringosc8[16].inv.y ;
 wire \tt_invring1.ringosc8[17].inv.y ;
 wire \tt_invring1.ringosc8[18].inv.y ;
 wire \tt_invring1.ringosc8[19].inv.y ;
 wire \tt_invring1.ringosc8[1].inv.y ;
 wire \tt_invring1.ringosc8[20].inv.y ;
 wire \tt_invring1.ringosc8[21].inv.y ;
 wire \tt_invring1.ringosc8[22].inv.y ;
 wire \tt_invring1.ringosc8[23].inv.y ;
 wire \tt_invring1.ringosc8[24].inv.y ;
 wire \tt_invring1.ringosc8[25].inv.y ;
 wire \tt_invring1.ringosc8[26].inv.y ;
 wire \tt_invring1.ringosc8[27].inv.y ;
 wire \tt_invring1.ringosc8[28].inv.y ;
 wire \tt_invring1.ringosc8[29].inv.y ;
 wire \tt_invring1.ringosc8[2].inv.y ;
 wire \tt_invring1.ringosc8[30].inv.y ;
 wire \tt_invring1.ringosc8[31].inv.y ;
 wire \tt_invring1.ringosc8[32].inv.y ;
 wire \tt_invring1.ringosc8[33].inv.y ;
 wire \tt_invring1.ringosc8[34].inv.y ;
 wire \tt_invring1.ringosc8[35].inv.y ;
 wire \tt_invring1.ringosc8[36].inv.y ;
 wire \tt_invring1.ringosc8[37].inv.y ;
 wire \tt_invring1.ringosc8[38].inv.y ;
 wire \tt_invring1.ringosc8[39].inv.y ;
 wire \tt_invring1.ringosc8[3].inv.y ;
 wire \tt_invring1.ringosc8[40].inv.y ;
 wire \tt_invring1.ringosc8[41].inv.y ;
 wire \tt_invring1.ringosc8[42].inv.y ;
 wire \tt_invring1.ringosc8[43].inv.y ;
 wire \tt_invring1.ringosc8[44].inv.y ;
 wire \tt_invring1.ringosc8[45].inv.y ;
 wire \tt_invring1.ringosc8[46].inv.y ;
 wire \tt_invring1.ringosc8[47].inv.y ;
 wire \tt_invring1.ringosc8[48].inv.y ;
 wire \tt_invring1.ringosc8[49].inv.y ;
 wire \tt_invring1.ringosc8[4].inv.y ;
 wire \tt_invring1.ringosc8[50].inv.y ;
 wire \tt_invring1.ringosc8[5].inv.y ;
 wire \tt_invring1.ringosc8[6].inv.y ;
 wire \tt_invring1.ringosc8[7].inv.y ;
 wire \tt_invring1.ringosc8[8].inv.y ;
 wire \tt_invring1.ringoutsam[0] ;
 wire \tt_invring1.ringoutsam[1] ;
 wire \tt_invring1.ringoutsam[2] ;
 wire \tt_invring1.ringoutsam[3] ;
 wire \tt_invring1.ringoutsam[4] ;
 wire \tt_invring1.ringoutsam[5] ;
 wire \tt_invring1.ringoutsam[6] ;
 wire \tt_invring1.ringoutsam[7] ;
 wire \tt_invring2.ringosc1[0].inv.a ;
 wire \tt_invring2.ringosc1[0].inv.y ;
 wire \tt_invring2.ringosc1[10].inv.a ;
 wire \tt_invring2.ringosc1[10].inv.y ;
 wire \tt_invring2.ringosc1[1].inv.y ;
 wire \tt_invring2.ringosc1[2].inv.y ;
 wire \tt_invring2.ringosc1[3].inv.y ;
 wire \tt_invring2.ringosc1[4].inv.y ;
 wire \tt_invring2.ringosc1[5].inv.y ;
 wire \tt_invring2.ringosc1[6].inv.y ;
 wire \tt_invring2.ringosc1[7].inv.y ;
 wire \tt_invring2.ringosc1[8].inv.y ;
 wire \tt_invring2.ringosc2[0].inv.a ;
 wire \tt_invring2.ringosc2[0].inv.y ;
 wire \tt_invring2.ringosc2[10].inv.a ;
 wire \tt_invring2.ringosc2[10].inv.y ;
 wire \tt_invring2.ringosc2[11].inv.y ;
 wire \tt_invring2.ringosc2[12].inv.y ;
 wire \tt_invring2.ringosc2[13].inv.y ;
 wire \tt_invring2.ringosc2[14].inv.y ;
 wire \tt_invring2.ringosc2[15].inv.y ;
 wire \tt_invring2.ringosc2[16].inv.y ;
 wire \tt_invring2.ringosc2[17].inv.y ;
 wire \tt_invring2.ringosc2[18].inv.y ;
 wire \tt_invring2.ringosc2[1].inv.y ;
 wire \tt_invring2.ringosc2[2].inv.y ;
 wire \tt_invring2.ringosc2[3].inv.y ;
 wire \tt_invring2.ringosc2[4].inv.y ;
 wire \tt_invring2.ringosc2[5].inv.y ;
 wire \tt_invring2.ringosc2[6].inv.y ;
 wire \tt_invring2.ringosc2[7].inv.y ;
 wire \tt_invring2.ringosc2[8].inv.y ;
 wire \tt_invring2.ringosc3[0].inv.a ;
 wire \tt_invring2.ringosc3[0].inv.y ;
 wire \tt_invring2.ringosc3[10].inv.a ;
 wire \tt_invring2.ringosc3[10].inv.y ;
 wire \tt_invring2.ringosc3[11].inv.y ;
 wire \tt_invring2.ringosc3[12].inv.y ;
 wire \tt_invring2.ringosc3[13].inv.y ;
 wire \tt_invring2.ringosc3[14].inv.y ;
 wire \tt_invring2.ringosc3[15].inv.y ;
 wire \tt_invring2.ringosc3[16].inv.y ;
 wire \tt_invring2.ringosc3[17].inv.y ;
 wire \tt_invring2.ringosc3[18].inv.y ;
 wire \tt_invring2.ringosc3[19].inv.y ;
 wire \tt_invring2.ringosc3[1].inv.y ;
 wire \tt_invring2.ringosc3[20].inv.y ;
 wire \tt_invring2.ringosc3[21].inv.y ;
 wire \tt_invring2.ringosc3[22].inv.y ;
 wire \tt_invring2.ringosc3[2].inv.y ;
 wire \tt_invring2.ringosc3[3].inv.y ;
 wire \tt_invring2.ringosc3[4].inv.y ;
 wire \tt_invring2.ringosc3[5].inv.y ;
 wire \tt_invring2.ringosc3[6].inv.y ;
 wire \tt_invring2.ringosc3[7].inv.y ;
 wire \tt_invring2.ringosc3[8].inv.y ;
 wire \tt_invring2.ringosc4[0].inv.a ;
 wire \tt_invring2.ringosc4[0].inv.y ;
 wire \tt_invring2.ringosc4[10].inv.a ;
 wire \tt_invring2.ringosc4[10].inv.y ;
 wire \tt_invring2.ringosc4[11].inv.y ;
 wire \tt_invring2.ringosc4[12].inv.y ;
 wire \tt_invring2.ringosc4[13].inv.y ;
 wire \tt_invring2.ringosc4[14].inv.y ;
 wire \tt_invring2.ringosc4[15].inv.y ;
 wire \tt_invring2.ringosc4[16].inv.y ;
 wire \tt_invring2.ringosc4[17].inv.y ;
 wire \tt_invring2.ringosc4[18].inv.y ;
 wire \tt_invring2.ringosc4[19].inv.y ;
 wire \tt_invring2.ringosc4[1].inv.y ;
 wire \tt_invring2.ringosc4[20].inv.y ;
 wire \tt_invring2.ringosc4[21].inv.y ;
 wire \tt_invring2.ringosc4[22].inv.y ;
 wire \tt_invring2.ringosc4[23].inv.y ;
 wire \tt_invring2.ringosc4[24].inv.y ;
 wire \tt_invring2.ringosc4[25].inv.y ;
 wire \tt_invring2.ringosc4[26].inv.y ;
 wire \tt_invring2.ringosc4[27].inv.y ;
 wire \tt_invring2.ringosc4[28].inv.y ;
 wire \tt_invring2.ringosc4[2].inv.y ;
 wire \tt_invring2.ringosc4[3].inv.y ;
 wire \tt_invring2.ringosc4[4].inv.y ;
 wire \tt_invring2.ringosc4[5].inv.y ;
 wire \tt_invring2.ringosc4[6].inv.y ;
 wire \tt_invring2.ringosc4[7].inv.y ;
 wire \tt_invring2.ringosc4[8].inv.y ;
 wire \tt_invring2.ringosc5[0].inv.a ;
 wire \tt_invring2.ringosc5[0].inv.y ;
 wire \tt_invring2.ringosc5[10].inv.a ;
 wire \tt_invring2.ringosc5[10].inv.y ;
 wire \tt_invring2.ringosc5[11].inv.y ;
 wire \tt_invring2.ringosc5[12].inv.y ;
 wire \tt_invring2.ringosc5[13].inv.y ;
 wire \tt_invring2.ringosc5[14].inv.y ;
 wire \tt_invring2.ringosc5[15].inv.y ;
 wire \tt_invring2.ringosc5[16].inv.y ;
 wire \tt_invring2.ringosc5[17].inv.y ;
 wire \tt_invring2.ringosc5[18].inv.y ;
 wire \tt_invring2.ringosc5[19].inv.y ;
 wire \tt_invring2.ringosc5[1].inv.y ;
 wire \tt_invring2.ringosc5[20].inv.y ;
 wire \tt_invring2.ringosc5[21].inv.y ;
 wire \tt_invring2.ringosc5[22].inv.y ;
 wire \tt_invring2.ringosc5[23].inv.y ;
 wire \tt_invring2.ringosc5[24].inv.y ;
 wire \tt_invring2.ringosc5[25].inv.y ;
 wire \tt_invring2.ringosc5[26].inv.y ;
 wire \tt_invring2.ringosc5[27].inv.y ;
 wire \tt_invring2.ringosc5[28].inv.y ;
 wire \tt_invring2.ringosc5[29].inv.y ;
 wire \tt_invring2.ringosc5[2].inv.y ;
 wire \tt_invring2.ringosc5[30].inv.y ;
 wire \tt_invring2.ringosc5[31].inv.y ;
 wire \tt_invring2.ringosc5[32].inv.y ;
 wire \tt_invring2.ringosc5[33].inv.y ;
 wire \tt_invring2.ringosc5[34].inv.y ;
 wire \tt_invring2.ringosc5[35].inv.y ;
 wire \tt_invring2.ringosc5[36].inv.y ;
 wire \tt_invring2.ringosc5[3].inv.y ;
 wire \tt_invring2.ringosc5[4].inv.y ;
 wire \tt_invring2.ringosc5[5].inv.y ;
 wire \tt_invring2.ringosc5[6].inv.y ;
 wire \tt_invring2.ringosc5[7].inv.y ;
 wire \tt_invring2.ringosc5[8].inv.y ;
 wire \tt_invring2.ringosc6[0].inv.a ;
 wire \tt_invring2.ringosc6[0].inv.y ;
 wire \tt_invring2.ringosc6[10].inv.a ;
 wire \tt_invring2.ringosc6[10].inv.y ;
 wire \tt_invring2.ringosc6[11].inv.y ;
 wire \tt_invring2.ringosc6[12].inv.y ;
 wire \tt_invring2.ringosc6[13].inv.y ;
 wire \tt_invring2.ringosc6[14].inv.y ;
 wire \tt_invring2.ringosc6[15].inv.y ;
 wire \tt_invring2.ringosc6[16].inv.y ;
 wire \tt_invring2.ringosc6[17].inv.y ;
 wire \tt_invring2.ringosc6[18].inv.y ;
 wire \tt_invring2.ringosc6[19].inv.y ;
 wire \tt_invring2.ringosc6[1].inv.y ;
 wire \tt_invring2.ringosc6[20].inv.y ;
 wire \tt_invring2.ringosc6[21].inv.y ;
 wire \tt_invring2.ringosc6[22].inv.y ;
 wire \tt_invring2.ringosc6[23].inv.y ;
 wire \tt_invring2.ringosc6[24].inv.y ;
 wire \tt_invring2.ringosc6[25].inv.y ;
 wire \tt_invring2.ringosc6[26].inv.y ;
 wire \tt_invring2.ringosc6[27].inv.y ;
 wire \tt_invring2.ringosc6[28].inv.y ;
 wire \tt_invring2.ringosc6[29].inv.y ;
 wire \tt_invring2.ringosc6[2].inv.y ;
 wire \tt_invring2.ringosc6[30].inv.y ;
 wire \tt_invring2.ringosc6[31].inv.y ;
 wire \tt_invring2.ringosc6[32].inv.y ;
 wire \tt_invring2.ringosc6[33].inv.y ;
 wire \tt_invring2.ringosc6[34].inv.y ;
 wire \tt_invring2.ringosc6[35].inv.y ;
 wire \tt_invring2.ringosc6[36].inv.y ;
 wire \tt_invring2.ringosc6[37].inv.y ;
 wire \tt_invring2.ringosc6[38].inv.y ;
 wire \tt_invring2.ringosc6[39].inv.y ;
 wire \tt_invring2.ringosc6[3].inv.y ;
 wire \tt_invring2.ringosc6[40].inv.y ;
 wire \tt_invring2.ringosc6[4].inv.y ;
 wire \tt_invring2.ringosc6[5].inv.y ;
 wire \tt_invring2.ringosc6[6].inv.y ;
 wire \tt_invring2.ringosc6[7].inv.y ;
 wire \tt_invring2.ringosc6[8].inv.y ;
 wire \tt_invring2.ringosc7[0].inv.a ;
 wire \tt_invring2.ringosc7[0].inv.y ;
 wire \tt_invring2.ringosc7[10].inv.a ;
 wire \tt_invring2.ringosc7[10].inv.y ;
 wire \tt_invring2.ringosc7[11].inv.y ;
 wire \tt_invring2.ringosc7[12].inv.y ;
 wire \tt_invring2.ringosc7[13].inv.y ;
 wire \tt_invring2.ringosc7[14].inv.y ;
 wire \tt_invring2.ringosc7[15].inv.y ;
 wire \tt_invring2.ringosc7[16].inv.y ;
 wire \tt_invring2.ringosc7[17].inv.y ;
 wire \tt_invring2.ringosc7[18].inv.y ;
 wire \tt_invring2.ringosc7[19].inv.y ;
 wire \tt_invring2.ringosc7[1].inv.y ;
 wire \tt_invring2.ringosc7[20].inv.y ;
 wire \tt_invring2.ringosc7[21].inv.y ;
 wire \tt_invring2.ringosc7[22].inv.y ;
 wire \tt_invring2.ringosc7[23].inv.y ;
 wire \tt_invring2.ringosc7[24].inv.y ;
 wire \tt_invring2.ringosc7[25].inv.y ;
 wire \tt_invring2.ringosc7[26].inv.y ;
 wire \tt_invring2.ringosc7[27].inv.y ;
 wire \tt_invring2.ringosc7[28].inv.y ;
 wire \tt_invring2.ringosc7[29].inv.y ;
 wire \tt_invring2.ringosc7[2].inv.y ;
 wire \tt_invring2.ringosc7[30].inv.y ;
 wire \tt_invring2.ringosc7[31].inv.y ;
 wire \tt_invring2.ringosc7[32].inv.y ;
 wire \tt_invring2.ringosc7[33].inv.y ;
 wire \tt_invring2.ringosc7[34].inv.y ;
 wire \tt_invring2.ringosc7[35].inv.y ;
 wire \tt_invring2.ringosc7[36].inv.y ;
 wire \tt_invring2.ringosc7[37].inv.y ;
 wire \tt_invring2.ringosc7[38].inv.y ;
 wire \tt_invring2.ringosc7[39].inv.y ;
 wire \tt_invring2.ringosc7[3].inv.y ;
 wire \tt_invring2.ringosc7[40].inv.y ;
 wire \tt_invring2.ringosc7[41].inv.y ;
 wire \tt_invring2.ringosc7[42].inv.y ;
 wire \tt_invring2.ringosc7[43].inv.y ;
 wire \tt_invring2.ringosc7[44].inv.y ;
 wire \tt_invring2.ringosc7[45].inv.y ;
 wire \tt_invring2.ringosc7[46].inv.y ;
 wire \tt_invring2.ringosc7[4].inv.y ;
 wire \tt_invring2.ringosc7[5].inv.y ;
 wire \tt_invring2.ringosc7[6].inv.y ;
 wire \tt_invring2.ringosc7[7].inv.y ;
 wire \tt_invring2.ringosc7[8].inv.y ;
 wire \tt_invring2.ringosc8[0].inv.a ;
 wire \tt_invring2.ringosc8[0].inv.y ;
 wire \tt_invring2.ringosc8[10].inv.a ;
 wire \tt_invring2.ringosc8[10].inv.y ;
 wire \tt_invring2.ringosc8[11].inv.y ;
 wire \tt_invring2.ringosc8[12].inv.y ;
 wire \tt_invring2.ringosc8[13].inv.y ;
 wire \tt_invring2.ringosc8[14].inv.y ;
 wire \tt_invring2.ringosc8[15].inv.y ;
 wire \tt_invring2.ringosc8[16].inv.y ;
 wire \tt_invring2.ringosc8[17].inv.y ;
 wire \tt_invring2.ringosc8[18].inv.y ;
 wire \tt_invring2.ringosc8[19].inv.y ;
 wire \tt_invring2.ringosc8[1].inv.y ;
 wire \tt_invring2.ringosc8[20].inv.y ;
 wire \tt_invring2.ringosc8[21].inv.y ;
 wire \tt_invring2.ringosc8[22].inv.y ;
 wire \tt_invring2.ringosc8[23].inv.y ;
 wire \tt_invring2.ringosc8[24].inv.y ;
 wire \tt_invring2.ringosc8[25].inv.y ;
 wire \tt_invring2.ringosc8[26].inv.y ;
 wire \tt_invring2.ringosc8[27].inv.y ;
 wire \tt_invring2.ringosc8[28].inv.y ;
 wire \tt_invring2.ringosc8[29].inv.y ;
 wire \tt_invring2.ringosc8[2].inv.y ;
 wire \tt_invring2.ringosc8[30].inv.y ;
 wire \tt_invring2.ringosc8[31].inv.y ;
 wire \tt_invring2.ringosc8[32].inv.y ;
 wire \tt_invring2.ringosc8[33].inv.y ;
 wire \tt_invring2.ringosc8[34].inv.y ;
 wire \tt_invring2.ringosc8[35].inv.y ;
 wire \tt_invring2.ringosc8[36].inv.y ;
 wire \tt_invring2.ringosc8[37].inv.y ;
 wire \tt_invring2.ringosc8[38].inv.y ;
 wire \tt_invring2.ringosc8[39].inv.y ;
 wire \tt_invring2.ringosc8[3].inv.y ;
 wire \tt_invring2.ringosc8[40].inv.y ;
 wire \tt_invring2.ringosc8[41].inv.y ;
 wire \tt_invring2.ringosc8[42].inv.y ;
 wire \tt_invring2.ringosc8[43].inv.y ;
 wire \tt_invring2.ringosc8[44].inv.y ;
 wire \tt_invring2.ringosc8[45].inv.y ;
 wire \tt_invring2.ringosc8[46].inv.y ;
 wire \tt_invring2.ringosc8[47].inv.y ;
 wire \tt_invring2.ringosc8[48].inv.y ;
 wire \tt_invring2.ringosc8[49].inv.y ;
 wire \tt_invring2.ringosc8[4].inv.y ;
 wire \tt_invring2.ringosc8[50].inv.y ;
 wire \tt_invring2.ringosc8[5].inv.y ;
 wire \tt_invring2.ringosc8[6].inv.y ;
 wire \tt_invring2.ringosc8[7].inv.y ;
 wire \tt_invring2.ringosc8[8].inv.y ;
 wire \tt_invring2.ringoutsam[0] ;
 wire \tt_invring2.ringoutsam[1] ;
 wire \tt_invring2.ringoutsam[2] ;
 wire \tt_invring2.ringoutsam[3] ;
 wire \tt_invring2.ringoutsam[4] ;
 wire \tt_invring2.ringoutsam[5] ;
 wire \tt_invring2.ringoutsam[6] ;
 wire \tt_invring2.ringoutsam[7] ;
 wire \tt_process.bitsadjacent[0] ;
 wire \tt_process.bitsadjacent[1] ;
 wire \tt_process.bitsadjacent[2] ;
 wire \tt_process.bitsgroup[0] ;
 wire \tt_process.bitsgroup[1] ;
 wire \tt_process.clk_half ;
 wire \tt_process.num ;
 wire \tt_process.tt_13n.connection[0] ;
 wire \tt_process.tt_13n.connection[10] ;
 wire \tt_process.tt_13n.connection[11] ;
 wire \tt_process.tt_13n.connection[12] ;
 wire \tt_process.tt_13n.connection[13] ;
 wire \tt_process.tt_13n.connection[1] ;
 wire \tt_process.tt_13n.connection[2] ;
 wire \tt_process.tt_13n.connection[3] ;
 wire \tt_process.tt_13n.connection[4] ;
 wire \tt_process.tt_13n.connection[5] ;
 wire \tt_process.tt_13n.connection[6] ;
 wire \tt_process.tt_13n.connection[7] ;
 wire \tt_process.tt_13n.connection[8] ;
 wire \tt_process.tt_13n.connection[9] ;
 wire \tt_samplekey.bitsadjacent[0] ;
 wire \tt_samplekey.bitsadjacent[1] ;
 wire \tt_samplekey.bitsadjacent[2] ;
 wire \tt_samplekey.bitsadjacent[3] ;
 wire \tt_samplekey.num ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;

 sky130_fd_sc_hd__and2_1 _138_ (.A(net41),
    .B(\tt_invring1.ringosc5[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc5[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _139_ (.A(net42),
    .B(\tt_invring1.ringosc4[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc4[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _140_ (.A(net42),
    .B(\tt_invring1.ringosc3[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc3[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _141_ (.A(net42),
    .B(\tt_invring1.ringosc2[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc2[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _142_ (.A(net42),
    .B(\tt_invring1.ringosc1[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc1[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _143_ (.A(net41),
    .B(\tt_invring2.ringosc8[50].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc8[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _144_ (.A(net41),
    .B(\tt_invring2.ringosc7[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc7[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _145_ (.A(net41),
    .B(\tt_invring2.ringosc6[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc6[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _146_ (.A(net41),
    .B(\tt_invring2.ringosc5[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc5[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _147_ (.A(net41),
    .B(\tt_invring2.ringosc4[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc4[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _148_ (.A(net41),
    .B(\tt_invring2.ringosc3[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc3[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _149_ (.A(net42),
    .B(\tt_invring2.ringosc2[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc2[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _150_ (.A(net42),
    .B(\tt_invring2.ringosc1[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring2.ringosc1[0].inv.a ));
 sky130_fd_sc_hd__nand2b_1 _151_ (.A_N(net92),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_007_));
 sky130_fd_sc_hd__and2_1 _152_ (.A(net46),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__and2_1 _153_ (.A(net46),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__and2_1 _154_ (.A(net46),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__and2_1 _155_ (.A(net44),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__and2_1 _156_ (.A(net47),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _157_ (.A(net44),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _158_ (.A(net45),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _159_ (.A(net44),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _160_ (.A(net44),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _161_ (.A(net44),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _162_ (.A(net46),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__and2_1 _163_ (.A(net46),
    .B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _164_ (.A(net46),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _165_ (.A(net46),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__and2_1 _166_ (.A(net47),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _167_ (.A(net49),
    .B(\tt_invring1.ringosc1[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _168_ (.A(net49),
    .B(\tt_invring1.ringosc2[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _169_ (.A(net49),
    .B(\tt_invring1.ringosc3[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__and2_1 _170_ (.A(net49),
    .B(\tt_invring1.ringosc4[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _171_ (.A(net43),
    .B(\tt_invring1.ringosc5[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__and2_1 _172_ (.A(net44),
    .B(\tt_invring1.ringosc6[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__and2_1 _173_ (.A(net46),
    .B(\tt_invring1.ringosc7[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__and2_1 _174_ (.A(net46),
    .B(\tt_invring1.ringosc8[50].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _175_ (.A(net48),
    .B(\tt_invring2.ringosc1[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__and2_1 _176_ (.A(net48),
    .B(\tt_invring2.ringosc2[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _177_ (.A(net43),
    .B(\tt_invring2.ringosc3[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _178_ (.A(net44),
    .B(\tt_invring2.ringosc4[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _179_ (.A(net44),
    .B(\tt_invring2.ringosc5[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _180_ (.A(net43),
    .B(\tt_invring2.ringosc6[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _181_ (.A(net44),
    .B(\tt_invring2.ringosc7[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__and2_1 _182_ (.A(net44),
    .B(\tt_invring2.ringosc8[50].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net48),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _184_ (.A(net48),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _185_ (.A(net48),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__and2_1 _186_ (.A(net45),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net45),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _188_ (.A(net45),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _189_ (.A(net45),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__and2_1 _190_ (.A(net47),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__and2_1 _191_ (.A(net47),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _192_ (.A(net49),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _193_ (.A(net49),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__and2_1 _194_ (.A(net49),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__and2_1 _195_ (.A(net49),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__and2_1 _196_ (.A(net48),
    .B(\tt_samplekey.num ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__and2_1 _197_ (.A(\tt_samplekey.bitsadjacent[0] ),
    .B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__and2_1 _198_ (.A(net9),
    .B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__and2_1 _199_ (.A(net8),
    .B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _200_ (.A(\tt_16bitran.connection[15] ),
    .B(\tt_16bitran.connection[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_135_));
 sky130_fd_sc_hd__xor2_1 _201_ (.A(\tt_16bitran.connection[13] ),
    .B(\tt_16bitran.connection[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__xnor2_1 _202_ (.A(_135_),
    .B(_136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_137_));
 sky130_fd_sc_hd__mux2_1 _203_ (.A0(net92),
    .A1(_137_),
    .S(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _204_ (.A0(\tt_process.tt_13n.connection[0] ),
    .A1(net66),
    .S(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__and2b_1 _205_ (.A_N(net91),
    .B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(\tt_samplekey.bitsadjacent[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(\tt_samplekey.bitsadjacent[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(\tt_process.bitsgroup[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_062_));
 sky130_fd_sc_hd__xnor2_1 _210_ (.A(\tt_invring1.ringoutsam[1] ),
    .B(\tt_invring1.ringoutsam[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_063_));
 sky130_fd_sc_hd__xor2_1 _211_ (.A(\tt_invring1.ringoutsam[2] ),
    .B(\tt_invring1.ringoutsam[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_064_));
 sky130_fd_sc_hd__xnor2_1 _212_ (.A(_063_),
    .B(_064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_065_));
 sky130_fd_sc_hd__xnor2_1 _213_ (.A(\tt_invring1.ringoutsam[6] ),
    .B(\tt_invring1.ringoutsam[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_066_));
 sky130_fd_sc_hd__xor2_1 _214_ (.A(\tt_invring1.ringoutsam[4] ),
    .B(\tt_invring1.ringoutsam[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(_066_),
    .B(_067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_068_));
 sky130_fd_sc_hd__a21oi_1 _216_ (.A1(net3),
    .A2(_065_),
    .B1(_068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_069_));
 sky130_fd_sc_hd__a31o_1 _217_ (.A1(net3),
    .A2(_065_),
    .A3(_068_),
    .B1(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(\tt_invring2.ringoutsam[6] ),
    .B(\tt_invring2.ringoutsam[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_071_));
 sky130_fd_sc_hd__xor2_1 _219_ (.A(\tt_invring2.ringoutsam[4] ),
    .B(\tt_invring2.ringoutsam[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_072_));
 sky130_fd_sc_hd__xnor2_1 _220_ (.A(_071_),
    .B(_072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_073_));
 sky130_fd_sc_hd__xor2_1 _221_ (.A(\tt_invring2.ringoutsam[2] ),
    .B(\tt_invring2.ringoutsam[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_074_));
 sky130_fd_sc_hd__xnor2_1 _222_ (.A(\tt_invring2.ringoutsam[1] ),
    .B(\tt_invring2.ringoutsam[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_075_));
 sky130_fd_sc_hd__xnor2_1 _223_ (.A(_074_),
    .B(_075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_076_));
 sky130_fd_sc_hd__a21oi_1 _224_ (.A1(net3),
    .A2(_076_),
    .B1(_073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_077_));
 sky130_fd_sc_hd__a31o_1 _225_ (.A1(net3),
    .A2(_073_),
    .A3(_076_),
    .B1(_059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__o22ai_1 _226_ (.A1(_069_),
    .A2(_070_),
    .B1(_077_),
    .B2(_078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_process.num ));
 sky130_fd_sc_hd__nand2_1 _227_ (.A(net9),
    .B(\tt_samplekey.bitsadjacent[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_079_));
 sky130_fd_sc_hd__a21o_1 _228_ (.A1(\tt_samplekey.bitsadjacent[2] ),
    .A2(_079_),
    .B1(\tt_samplekey.bitsadjacent[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_080_));
 sky130_fd_sc_hd__o21ba_1 _229_ (.A1(net9),
    .A2(_060_),
    .B1_N(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__nand2_1 _230_ (.A(\tt_samplekey.bitsadjacent[2] ),
    .B(\tt_samplekey.bitsadjacent[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_082_));
 sky130_fd_sc_hd__o32a_1 _231_ (.A1(\tt_samplekey.bitsadjacent[1] ),
    .A2(\tt_samplekey.bitsadjacent[0] ),
    .A3(_082_),
    .B1(_081_),
    .B2(_080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_000_));
 sky130_fd_sc_hd__o31a_1 _232_ (.A1(\tt_samplekey.bitsadjacent[1] ),
    .A2(_060_),
    .A3(_082_),
    .B1(_080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__nor2_1 _233_ (.A(net9),
    .B(\tt_samplekey.bitsadjacent[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _234_ (.A(net8),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_084_));
 sky130_fd_sc_hd__o22ai_1 _235_ (.A1(\tt_samplekey.bitsadjacent[0] ),
    .A2(_083_),
    .B1(_084_),
    .B2(_061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_1 _236_ (.A(net8),
    .B(_061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_085_));
 sky130_fd_sc_hd__mux2_1 _237_ (.A0(net8),
    .A1(_085_),
    .S(_060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(_083_),
    .A1(net9),
    .S(_086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_087_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(_087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _240_ (.A(net8),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_088_));
 sky130_fd_sc_hd__o21a_1 _241_ (.A1(\tt_samplekey.bitsadjacent[0] ),
    .A2(_085_),
    .B1(_088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_089_));
 sky130_fd_sc_hd__a21o_1 _242_ (.A1(net8),
    .A2(_061_),
    .B1(_089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__and2_1 _243_ (.A(net8),
    .B(_083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_090_));
 sky130_fd_sc_hd__a21oi_1 _244_ (.A1(net9),
    .A2(\tt_samplekey.bitsadjacent[3] ),
    .B1(_090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_091_));
 sky130_fd_sc_hd__o21ai_1 _245_ (.A1(net8),
    .A2(_083_),
    .B1(_060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_092_));
 sky130_fd_sc_hd__o22a_1 _246_ (.A1(_060_),
    .A2(_091_),
    .B1(_092_),
    .B2(_090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__or4b_1 _247_ (.A(_060_),
    .B(_061_),
    .C(_084_),
    .D_N(_088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_093_));
 sky130_fd_sc_hd__o31a_1 _248_ (.A1(net9),
    .A2(\tt_samplekey.bitsadjacent[3] ),
    .A3(_086_),
    .B1(_093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _249_ (.A0(\tt_finalprocess.genblk1[7].multblock.multblockout ),
    .A1(\tt_finalprocess.genblk1[3].multblock.multblockout ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_094_));
 sky130_fd_sc_hd__and2_2 _250_ (.A(net43),
    .B(_094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_095_));
 sky130_fd_sc_hd__nand2_1 _251_ (.A(net43),
    .B(_094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_096_));
 sky130_fd_sc_hd__mux2_1 _252_ (.A0(\tt_finalprocess.genblk1[6].multblock.multblockout ),
    .A1(\tt_finalprocess.genblk1[2].multblock.multblockout ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_097_));
 sky130_fd_sc_hd__and2_1 _253_ (.A(net43),
    .B(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_098_));
 sky130_fd_sc_hd__nand2_1 _254_ (.A(net43),
    .B(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_099_));
 sky130_fd_sc_hd__mux2_1 _255_ (.A0(\tt_finalprocess.genblk1[5].multblock.multblockout ),
    .A1(\tt_finalprocess.genblk1[1].multblock.multblockout ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_100_));
 sky130_fd_sc_hd__and2_1 _256_ (.A(net43),
    .B(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_101_));
 sky130_fd_sc_hd__nand2_2 _257_ (.A(net43),
    .B(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_102_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\tt_finalprocess.genblk1[4].multblock.multblockout ),
    .A1(\tt_finalprocess.genblk1[0].multblock.multblockout ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_103_));
 sky130_fd_sc_hd__nand2_1 _259_ (.A(net43),
    .B(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_104_));
 sky130_fd_sc_hd__and3_1 _260_ (.A(_098_),
    .B(_102_),
    .C(_104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_105_));
 sky130_fd_sc_hd__nor2_2 _261_ (.A(_101_),
    .B(_104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _262_ (.A(_098_),
    .B(_106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_107_));
 sky130_fd_sc_hd__and3_1 _263_ (.A(net1),
    .B(_100_),
    .C(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(_099_),
    .B(_108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_109_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(_095_),
    .B(_109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_110_));
 sky130_fd_sc_hd__o2bb2a_4 _266_ (.A1_N(_095_),
    .A2_N(_105_),
    .B1(_107_),
    .B2(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__and3_1 _267_ (.A(net1),
    .B(_097_),
    .C(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_111_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(_111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_112_));
 sky130_fd_sc_hd__o31a_4 _269_ (.A1(_096_),
    .A2(_101_),
    .A3(_112_),
    .B1(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__o21a_1 _270_ (.A1(_102_),
    .A2(_103_),
    .B1(_096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__nor2_1 _271_ (.A(_096_),
    .B(_098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_114_));
 sky130_fd_sc_hd__a21oi_4 _272_ (.A1(_106_),
    .A2(_114_),
    .B1(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uio_out[2]));
 sky130_fd_sc_hd__or3_1 _273_ (.A(_095_),
    .B(_101_),
    .C(_111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__or4_1 _274_ (.A(_096_),
    .B(_098_),
    .C(_102_),
    .D(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__o211a_4 _275_ (.A1(_102_),
    .A2(_112_),
    .B1(_115_),
    .C1(_116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__a21oi_1 _276_ (.A1(_099_),
    .A2(_104_),
    .B1(_095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_117_));
 sky130_fd_sc_hd__or3_4 _277_ (.A(_106_),
    .B(_114_),
    .C(_117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__o21ai_1 _278_ (.A1(_098_),
    .A2(_108_),
    .B1(_095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_118_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(_102_),
    .A2(_104_),
    .B1(_109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_119_));
 sky130_fd_sc_hd__o32a_4 _280_ (.A1(_095_),
    .A2(_105_),
    .A3(_119_),
    .B1(_118_),
    .B2(_106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__nor2_1 _281_ (.A(_099_),
    .B(_106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_120_));
 sky130_fd_sc_hd__o21a_2 _282_ (.A1(_118_),
    .A2(_120_),
    .B1(_115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(\tt_process.tt_13n.connection[10] ),
    .B(\tt_process.tt_13n.connection[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_121_));
 sky130_fd_sc_hd__xor2_1 _284_ (.A(\tt_process.tt_13n.connection[3] ),
    .B(\tt_process.tt_13n.connection[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__xnor2_1 _285_ (.A(\tt_process.tt_13n.connection[5] ),
    .B(_122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_123_));
 sky130_fd_sc_hd__xnor2_1 _286_ (.A(_121_),
    .B(_123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_124_));
 sky130_fd_sc_hd__xor2_1 _287_ (.A(\tt_process.tt_13n.connection[7] ),
    .B(\tt_process.tt_13n.connection[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__xor2_1 _288_ (.A(\tt_process.tt_13n.connection[2] ),
    .B(\tt_process.tt_13n.connection[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__xnor2_1 _289_ (.A(_125_),
    .B(_126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_127_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(\tt_process.tt_13n.connection[12] ),
    .B(\tt_process.tt_13n.connection[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_128_));
 sky130_fd_sc_hd__xor2_1 _291_ (.A(\tt_process.tt_13n.connection[6] ),
    .B(\tt_process.tt_13n.connection[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__xnor2_1 _292_ (.A(_128_),
    .B(_129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_130_));
 sky130_fd_sc_hd__xnor2_1 _293_ (.A(_127_),
    .B(_130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_131_));
 sky130_fd_sc_hd__nand2_1 _294_ (.A(_124_),
    .B(_131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_132_));
 sky130_fd_sc_hd__o22a_1 _295_ (.A1(\tt_process.bitsgroup[0] ),
    .A2(_062_),
    .B1(_124_),
    .B2(_131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__a22o_1 _296_ (.A1(\tt_process.bitsgroup[0] ),
    .A2(_062_),
    .B1(_132_),
    .B2(_133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__xnor2_2 _297_ (.A(\tt_16bitran.connection[0] ),
    .B(_134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_samplekey.num ));
 sky130_fd_sc_hd__and2_1 _298_ (.A(\tt_invring1.ringosc8[50].inv.y ),
    .B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc8[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _299_ (.A(net41),
    .B(\tt_invring1.ringosc7[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc7[0].inv.a ));
 sky130_fd_sc_hd__and2_1 _300_ (.A(net41),
    .B(\tt_invring1.ringosc6[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_invring1.ringosc6[0].inv.a ));
 sky130_fd_sc_hd__dfxtp_1 _301_ (.CLK(clknet_2_1__leaf_clk),
    .D(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[1] ));
 sky130_fd_sc_hd__dfxtp_1 _302_ (.CLK(clknet_2_1__leaf_clk),
    .D(_008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[2] ));
 sky130_fd_sc_hd__dfxtp_1 _303_ (.CLK(clknet_2_1__leaf_clk),
    .D(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[3] ));
 sky130_fd_sc_hd__dfxtp_1 _304_ (.CLK(clknet_2_1__leaf_clk),
    .D(_010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[4] ));
 sky130_fd_sc_hd__dfxtp_1 _305_ (.CLK(clknet_2_0__leaf_clk),
    .D(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[5] ));
 sky130_fd_sc_hd__dfxtp_1 _306_ (.CLK(clknet_2_0__leaf_clk),
    .D(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[6] ));
 sky130_fd_sc_hd__dfxtp_1 _307_ (.CLK(clknet_2_0__leaf_clk),
    .D(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[7] ));
 sky130_fd_sc_hd__dfxtp_1 _308_ (.CLK(clknet_2_1__leaf_clk),
    .D(_014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[8] ));
 sky130_fd_sc_hd__dfxtp_1 _309_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[9] ));
 sky130_fd_sc_hd__dfxtp_1 _310_ (.CLK(clknet_2_0__leaf_clk),
    .D(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[10] ));
 sky130_fd_sc_hd__dfxtp_1 _311_ (.CLK(clknet_2_0__leaf_clk),
    .D(_017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[11] ));
 sky130_fd_sc_hd__dfxtp_1 _312_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[12] ));
 sky130_fd_sc_hd__dfxtp_1 _313_ (.CLK(clknet_2_1__leaf_clk),
    .D(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[13] ));
 sky130_fd_sc_hd__dfxtp_1 _314_ (.CLK(clknet_2_1__leaf_clk),
    .D(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[14] ));
 sky130_fd_sc_hd__dfxtp_1 _315_ (.CLK(clknet_2_1__leaf_clk),
    .D(_021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[15] ));
 sky130_fd_sc_hd__dfxtp_1 _316_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[16] ));
 sky130_fd_sc_hd__dfxtp_1 _317_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[0] ));
 sky130_fd_sc_hd__dfxtp_1 _318_ (.CLK(clknet_2_3__leaf_clk),
    .D(_024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[1] ));
 sky130_fd_sc_hd__dfxtp_1 _319_ (.CLK(clknet_2_3__leaf_clk),
    .D(_025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[2] ));
 sky130_fd_sc_hd__dfxtp_1 _320_ (.CLK(clknet_2_3__leaf_clk),
    .D(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[3] ));
 sky130_fd_sc_hd__dfxtp_1 _321_ (.CLK(clknet_2_0__leaf_clk),
    .D(_027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[4] ));
 sky130_fd_sc_hd__dfxtp_1 _322_ (.CLK(clknet_2_0__leaf_clk),
    .D(_028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[5] ));
 sky130_fd_sc_hd__dfxtp_1 _323_ (.CLK(clknet_2_1__leaf_clk),
    .D(_029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[6] ));
 sky130_fd_sc_hd__dfxtp_1 _324_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring1.ringoutsam[7] ));
 sky130_fd_sc_hd__dfxtp_1 _325_ (.CLK(clknet_2_2__leaf_clk),
    .D(_031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[0] ));
 sky130_fd_sc_hd__dfxtp_1 _326_ (.CLK(clknet_2_2__leaf_clk),
    .D(_032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[1] ));
 sky130_fd_sc_hd__dfxtp_1 _327_ (.CLK(clknet_2_0__leaf_clk),
    .D(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[2] ));
 sky130_fd_sc_hd__dfxtp_1 _328_ (.CLK(clknet_2_0__leaf_clk),
    .D(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[3] ));
 sky130_fd_sc_hd__dfxtp_1 _329_ (.CLK(clknet_2_0__leaf_clk),
    .D(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[4] ));
 sky130_fd_sc_hd__dfxtp_1 _330_ (.CLK(clknet_2_0__leaf_clk),
    .D(_036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[5] ));
 sky130_fd_sc_hd__dfxtp_1 _331_ (.CLK(clknet_2_0__leaf_clk),
    .D(_037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[6] ));
 sky130_fd_sc_hd__dfxtp_1 _332_ (.CLK(clknet_2_1__leaf_clk),
    .D(_038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_invring2.ringoutsam[7] ));
 sky130_fd_sc_hd__dfxtp_1 _333_ (.CLK(\tt_process.clk_half ),
    .D(\tt_process.bitsadjacent[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.bitsgroup[0] ));
 sky130_fd_sc_hd__dfxtp_1 _334_ (.CLK(\tt_process.clk_half ),
    .D(\tt_process.bitsadjacent[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.bitsgroup[1] ));
 sky130_fd_sc_hd__dfxtp_1 _335_ (.CLK(clknet_2_3__leaf_clk),
    .D(\tt_process.num ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.bitsadjacent[0] ));
 sky130_fd_sc_hd__dfxtp_1 _336_ (.CLK(clknet_2_3__leaf_clk),
    .D(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.bitsadjacent[1] ));
 sky130_fd_sc_hd__dfxtp_1 _337_ (.CLK(clknet_2_2__leaf_clk),
    .D(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.bitsadjacent[2] ));
 sky130_fd_sc_hd__dfxtp_2 _338_ (.CLK(net40),
    .D(_000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_2 _339_ (.CLK(net40),
    .D(_001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_2 _340_ (.CLK(net40),
    .D(_002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _341_ (.CLK(net40),
    .D(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _342_ (.CLK(net40),
    .D(_004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _343_ (.CLK(net40),
    .D(_005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _344_ (.CLK(net40),
    .D(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_1 _345_ (.CLK(clknet_2_2__leaf_clk),
    .D(_039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[1] ));
 sky130_fd_sc_hd__dfxtp_1 _346_ (.CLK(clknet_2_2__leaf_clk),
    .D(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[2] ));
 sky130_fd_sc_hd__dfxtp_1 _347_ (.CLK(clknet_2_2__leaf_clk),
    .D(_041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[3] ));
 sky130_fd_sc_hd__dfxtp_1 _348_ (.CLK(clknet_2_0__leaf_clk),
    .D(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[4] ));
 sky130_fd_sc_hd__dfxtp_1 _349_ (.CLK(clknet_2_0__leaf_clk),
    .D(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[5] ));
 sky130_fd_sc_hd__dfxtp_1 _350_ (.CLK(clknet_2_2__leaf_clk),
    .D(_044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[6] ));
 sky130_fd_sc_hd__dfxtp_1 _351_ (.CLK(clknet_2_0__leaf_clk),
    .D(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[7] ));
 sky130_fd_sc_hd__dfxtp_1 _352_ (.CLK(clknet_2_1__leaf_clk),
    .D(_046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[8] ));
 sky130_fd_sc_hd__dfxtp_1 _353_ (.CLK(clknet_2_1__leaf_clk),
    .D(_047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[9] ));
 sky130_fd_sc_hd__dfxtp_1 _354_ (.CLK(clknet_2_3__leaf_clk),
    .D(_048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[10] ));
 sky130_fd_sc_hd__dfxtp_1 _355_ (.CLK(clknet_2_3__leaf_clk),
    .D(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[11] ));
 sky130_fd_sc_hd__dfxtp_1 _356_ (.CLK(clknet_2_3__leaf_clk),
    .D(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[12] ));
 sky130_fd_sc_hd__dfxtp_1 _357_ (.CLK(clknet_2_1__leaf_clk),
    .D(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[13] ));
 sky130_fd_sc_hd__dfxtp_1 _358_ (.CLK(net5),
    .D(\tt_samplekey.bitsadjacent[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.key ));
 sky130_fd_sc_hd__dfxtp_1 _359_ (.CLK(net40),
    .D(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.key ));
 sky130_fd_sc_hd__dfxtp_1 _360_ (.CLK(net40),
    .D(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.key ));
 sky130_fd_sc_hd__dfxtp_1 _361_ (.CLK(net40),
    .D(\tt_samplekey.bitsadjacent[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.key ));
 sky130_fd_sc_hd__dfxtp_1 _362_ (.CLK(clknet_2_2__leaf_clk),
    .D(_052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_samplekey.bitsadjacent[0] ));
 sky130_fd_sc_hd__dfxtp_1 _363_ (.CLK(clknet_2_2__leaf_clk),
    .D(_053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_samplekey.bitsadjacent[1] ));
 sky130_fd_sc_hd__dfxtp_1 _364_ (.CLK(clknet_2_2__leaf_clk),
    .D(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_samplekey.bitsadjacent[2] ));
 sky130_fd_sc_hd__dfxtp_2 _365_ (.CLK(clknet_2_3__leaf_clk),
    .D(_055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_samplekey.bitsadjacent[3] ));
 sky130_fd_sc_hd__dfxtp_1 _366_ (.CLK(clknet_2_1__leaf_clk),
    .D(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_16bitran.connection[0] ));
 sky130_fd_sc_hd__dfxtp_1 _367_ (.CLK(clknet_2_2__leaf_clk),
    .D(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.tt_13n.connection[0] ));
 sky130_fd_sc_hd__dfxtp_1 _368_ (.CLK(clknet_2_2__leaf_clk),
    .D(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tt_process.clk_half ));
 sky130_fd_sc_hd__buf_2 _369_ (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _370_ (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _371_ (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _372_ (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__buf_2 _373_ (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__buf_2 _374_ (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__buf_2 _375_ (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _376_ (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__clkbuf_4 _377_ (.A(\tt_samplekey.num ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__clkbuf_4 _378_ (.A(\tt_process.num ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net39),
    .A1(net39),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net39),
    .A1(net39),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.b ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.a ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.d ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.c ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.d ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.c ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.d ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[1].mult_22.c ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.d ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[2].mult_22.c ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.d ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.c ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.d ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[4].mult_22.c ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.d ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[5].mult_22.c ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.d ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.c ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.d ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[7].mult_22.c ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.d ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[0].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[0].multblock.genblk1[8].mult_22.c ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[0].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[0].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[0].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[0].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[0].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[0].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[0].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net36),
    .A1(net36),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net37),
    .A1(net37),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.b ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.a ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.d ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.c ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.d ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[0].mult_22.c ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.d ),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[1].mult_22.c ),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.d ),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[2].mult_22.c ),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.d ),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[3].mult_22.c ),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.d ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[4].mult_22.c ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.d ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[5].mult_22.c ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.d ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[6].mult_22.c ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.d ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[7].mult_22.c ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.d ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[1].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[1].multblock.genblk1[8].mult_22.c ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[1].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[1].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[1].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[1].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[1].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[1].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[1].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[1].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net36),
    .A1(net36),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net36),
    .A1(net36),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.b ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.a ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.d ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.c ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.d ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[0].mult_22.c ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.d ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[1].mult_22.c ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.d ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[2].mult_22.c ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.d ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[3].mult_22.c ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.d ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[4].mult_22.c ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.d ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[5].mult_22.c ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.d ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[6].mult_22.c ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.d ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[7].mult_22.c ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.d ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[2].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[2].multblock.genblk1[8].mult_22.c ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[2].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[2].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[2].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[2].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[2].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[2].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[2].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[2].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net39),
    .A1(net39),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net6),
    .A1(net6),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.b ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.a ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.d ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.c ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.d ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[0].mult_22.c ),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.d ),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[1].mult_22.c ),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.d ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[2].mult_22.c ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.d ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[3].mult_22.c ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.d ),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[4].mult_22.c ),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.d ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[5].mult_22.c ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.d ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[6].mult_22.c ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.d ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[7].mult_22.c ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.d ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[3].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[3].multblock.genblk1[8].mult_22.c ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[3].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[3].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[3].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[3].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[3].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[3].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[3].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[3].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net39),
    .A1(net39),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net39),
    .A1(net39),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.b ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.a ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.d ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.c ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.d ),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[0].mult_22.c ),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.d ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[1].mult_22.c ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.d ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[2].mult_22.c ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.d ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[3].mult_22.c ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.d ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[4].mult_22.c ),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.d ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[5].mult_22.c ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.d ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[6].mult_22.c ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.d ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[7].mult_22.c ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.d ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[4].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[4].multblock.genblk1[8].mult_22.c ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[4].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[4].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[4].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[4].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[4].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[4].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[4].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[4].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net38),
    .A1(net38),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net38),
    .A1(net38),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.b ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.a ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.d ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.c ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.d ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[0].mult_22.c ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.d ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[1].mult_22.c ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.d ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[2].mult_22.c ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.d ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[3].mult_22.c ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.d ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[4].mult_22.c ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.d ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[5].mult_22.c ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.d ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[6].mult_22.c ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.d ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[7].mult_22.c ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.d ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[5].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[5].multblock.genblk1[8].mult_22.c ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[5].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[5].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[5].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[5].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[5].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[5].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[5].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[5].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net36),
    .A1(net36),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net36),
    .A1(net36),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.b ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.a ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.d ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.c ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.d ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[0].mult_22.c ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.d ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[1].mult_22.c ),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.d ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[2].mult_22.c ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.d ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[3].mult_22.c ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.d ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[4].mult_22.c ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.d ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[5].mult_22.c ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.d ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[6].mult_22.c ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.d ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[7].mult_22.c ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.d ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[6].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[6].multblock.genblk1[8].mult_22.c ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[6].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[6].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[6].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[6].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[6].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[6].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[6].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[6].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.mult_1.cell0_I  (.A0(net37),
    .A1(net37),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.mult_2.cell0_I  (.A0(net37),
    .A1(net37),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.a ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.b ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.b ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.a ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.d ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.c ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.d ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[0].mult_22.c ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.d ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[1].mult_22.c ),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.d ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[2].mult_22.c ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.d ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[3].mult_22.c ),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.d ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[4].mult_22.c ),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.d ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[5].mult_22.c ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.d ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[6].mult_22.c ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.d ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.c ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[7].mult_22.c ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.d ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[9].mult_22.mult_1.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.c ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.d ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.a ));
 sky130_fd_sc_hd__mux2_1 \tt_finalprocess.genblk1[7].multblock.genblk1[9].mult_22.mult_2.cell0_I  (.A0(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.d ),
    .A1(\tt_finalprocess.genblk1[7].multblock.genblk1[8].mult_22.c ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tt_finalprocess.genblk1[7].multblock.genblk1[10].mult_22.b ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[7].multblock.nand_gate_2.nand_gate1.cell_nand  (.A(\tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.c ),
    .B(\tt_finalprocess.genblk1[7].multblock.nand_gate_2.B_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[7].multblock.multblockout ));
 sky130_fd_sc_hd__nand2_1 \tt_finalprocess.genblk1[7].multblock.nand_gate_2.nand_gate2.cell_nand  (.A(\tt_finalprocess.genblk1[7].multblock.multblockout ),
    .B(\tt_finalprocess.genblk1[7].multblock.genblk1[11].mult_22.d ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_finalprocess.genblk1[7].multblock.nand_gate_2.B_1 ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc1[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc1[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc1[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc2[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc2[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc2[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc3[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc3[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc3[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[23].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[24].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[25].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[26].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[27].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[28].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc4[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc4[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc4[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[23].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[24].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[25].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[26].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[27].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[28].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[29].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[30].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[31].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[32].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[33].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[34].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[35].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[36].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc5[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc5[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc5[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[23].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[24].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[25].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[26].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[27].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[28].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[29].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[30].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[31].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[32].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[33].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[34].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[35].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[36].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[37].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[38].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[39].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[40].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc6[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc6[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc6[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[23].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[24].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[25].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[26].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[27].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[28].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[29].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[30].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[31].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[32].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[33].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[34].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[35].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[36].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[37].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[38].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[39].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[40].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[41].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[41].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[42].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[41].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[42].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[43].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[42].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[43].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[44].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[43].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[44].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[45].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[44].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[45].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[46].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[45].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[46].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc7[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc7[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc7[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[0].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[10].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[11].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[12].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[13].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[14].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[15].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[16].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[17].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[18].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[19].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[1].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[20].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[21].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[22].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[23].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[24].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[25].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[26].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[27].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[28].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[29].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[2].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[30].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[31].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[32].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[33].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[34].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[35].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[36].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[37].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[38].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[39].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[3].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[40].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[41].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[41].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[42].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[41].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[42].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[43].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[42].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[43].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[44].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[43].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[44].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[45].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[44].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[45].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[46].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[45].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[46].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[47].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[47].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[48].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[47].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[48].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[49].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[48].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[49].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[4].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[50].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[49].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[50].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[5].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[6].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[7].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[8].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring1.ringosc8[9].inv.cnt_bit_I  (.A(\tt_invring1.ringosc8[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring1.ringosc8[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc1[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc1[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc1[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc2[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc2[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc2[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc3[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc3[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc3[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[23].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[24].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[25].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[26].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[27].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[28].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc4[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc4[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc4[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[23].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[24].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[25].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[26].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[27].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[28].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[29].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[30].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[31].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[32].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[33].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[34].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[35].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[36].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc5[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc5[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc5[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[23].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[24].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[25].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[26].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[27].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[28].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[29].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[30].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[31].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[32].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[33].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[34].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[35].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[36].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[37].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[38].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[39].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[40].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc6[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc6[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc6[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[23].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[24].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[25].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[26].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[27].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[28].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[29].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[30].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[31].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[32].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[33].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[34].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[35].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[36].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[37].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[38].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[39].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[40].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[41].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[41].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[42].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[41].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[42].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[43].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[42].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[43].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[44].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[43].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[44].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[45].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[44].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[45].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[46].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[45].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[46].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc7[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc7[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc7[10].inv.a ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[0].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[0].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[0].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[10].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[10].inv.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[10].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[11].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[10].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[11].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[12].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[11].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[12].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[13].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[12].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[13].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[14].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[13].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[14].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[15].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[14].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[15].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[16].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[15].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[16].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[17].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[16].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[17].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[18].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[17].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[18].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[19].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[18].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[19].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[1].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[0].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[1].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[20].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[19].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[20].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[21].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[20].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[21].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[22].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[21].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[22].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[23].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[22].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[23].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[24].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[23].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[24].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[25].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[24].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[25].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[26].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[25].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[26].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[27].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[26].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[27].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[28].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[27].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[28].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[29].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[28].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[29].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[2].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[1].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[2].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[30].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[29].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[30].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[31].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[30].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[31].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[32].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[31].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[32].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[33].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[32].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[33].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[34].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[33].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[34].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[35].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[34].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[35].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[36].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[35].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[36].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[37].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[36].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[37].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[38].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[37].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[38].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[39].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[38].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[39].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[3].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[2].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[3].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[40].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[39].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[40].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[41].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[40].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[41].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[42].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[41].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[42].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[43].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[42].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[43].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[44].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[43].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[44].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[45].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[44].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[45].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[46].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[45].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[46].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[47].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[46].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[47].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[48].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[47].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[48].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[49].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[48].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[49].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[4].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[3].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[4].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[50].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[49].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[50].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[5].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[4].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[5].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[6].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[5].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[6].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[7].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[6].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[7].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[8].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[7].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[8].inv.y ));
 sky130_fd_sc_hd__inv_2 \tt_invring2.ringosc8[9].inv.cnt_bit_I  (.A(\tt_invring2.ringosc8[8].inv.y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tt_invring2.ringosc8[10].inv.a ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 fanout8 (.A(\tt_samplekey.bitsadjacent[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_2 fanout9 (.A(\tt_samplekey.bitsadjacent[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[10].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout21 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout22 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[6].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[3].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(\tt_finalprocess.genblk1[0].multblock.genblk1[0].mult_22.key ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_1 fanout37 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_1 fanout38 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout42 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_1 fanout45 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_1 fanout47 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__conb_1 _369__51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net51));
 sky130_fd_sc_hd__conb_1 _370__52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net52));
 sky130_fd_sc_hd__conb_1 _371__53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net53));
 sky130_fd_sc_hd__conb_1 _372__54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net54));
 sky130_fd_sc_hd__conb_1 _373__55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net55));
 sky130_fd_sc_hd__conb_1 _374__56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net56));
 sky130_fd_sc_hd__conb_1 _375__57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net57));
 sky130_fd_sc_hd__conb_1 _376__58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net58));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\tt_process.bitsadjacent[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\tt_process.bitsadjacent[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\tt_16bitran.connection[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\tt_16bitran.connection[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\tt_16bitran.connection[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\tt_16bitran.connection[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\tt_16bitran.connection[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\tt_process.bitsadjacent[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\tt_16bitran.connection[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\tt_16bitran.connection[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\tt_16bitran.connection[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\tt_16bitran.connection[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\tt_16bitran.connection[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\tt_16bitran.connection[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\tt_16bitran.connection[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\tt_process.tt_13n.connection[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\tt_process.tt_13n.connection[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\tt_process.tt_13n.connection[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\tt_process.tt_13n.connection[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\tt_process.tt_13n.connection[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\tt_process.tt_13n.connection[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\tt_process.tt_13n.connection[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\tt_process.tt_13n.connection[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\tt_process.tt_13n.connection[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\tt_16bitran.connection[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\tt_process.tt_13n.connection[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\tt_process.tt_13n.connection[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\tt_16bitran.connection[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\tt_process.tt_13n.connection[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\tt_process.tt_13n.connection[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\tt_16bitran.connection[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\tt_process.clk_half ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\tt_16bitran.connection[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_295 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_200 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_308 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_147 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_217 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_268 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_166 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_222 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_234 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_159 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_159 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_171 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_208 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_220 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_232 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_190 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_106 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_194 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_55 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_129 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_66 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_284 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_84 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_247 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_217 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_136 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_256 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_213 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_13 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_167 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_145 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_210 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_16 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_32 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_107 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_210 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_271 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
