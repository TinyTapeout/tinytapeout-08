VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 1349.361206 ;
    ANTENNADIFFAREA 520.631958 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    USE POWER ;
    ANTENNAGATEAREA 853.044495 ;
    ANTENNADIFFAREA 1113.359375 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.725 211.225 14.895 211.415 ;
        RECT 18.405 211.225 18.575 211.415 ;
        RECT 23.925 211.225 24.095 211.415 ;
        RECT 25.765 211.225 25.935 211.415 ;
        RECT 31.285 211.225 31.455 211.415 ;
        RECT 36.805 211.225 36.975 211.415 ;
        RECT 38.645 211.225 38.815 211.415 ;
        RECT 44.165 211.225 44.335 211.415 ;
        RECT 49.685 211.225 49.855 211.415 ;
        RECT 51.525 211.225 51.695 211.415 ;
        RECT 57.045 211.225 57.215 211.415 ;
        RECT 62.565 211.225 62.735 211.415 ;
        RECT 64.405 211.225 64.575 211.415 ;
        RECT 69.925 211.225 70.095 211.415 ;
        RECT 75.445 211.225 75.615 211.415 ;
        RECT 77.285 211.225 77.455 211.415 ;
        RECT 82.805 211.225 82.975 211.415 ;
        RECT 88.325 211.225 88.495 211.415 ;
        RECT 90.165 211.225 90.335 211.415 ;
        RECT 95.685 211.225 95.855 211.415 ;
        RECT 101.205 211.225 101.375 211.415 ;
        RECT 103.045 211.225 103.215 211.415 ;
        RECT 108.565 211.225 108.735 211.415 ;
        RECT 114.085 211.225 114.255 211.415 ;
        RECT 115.060 211.275 115.180 211.385 ;
        RECT 120.525 211.225 120.695 211.415 ;
        RECT 126.045 211.225 126.215 211.415 ;
        RECT 127.425 211.225 127.595 211.415 ;
        RECT 14.585 210.415 15.955 211.225 ;
        RECT 15.965 210.415 18.715 211.225 ;
        RECT 18.725 210.415 24.235 211.225 ;
        RECT 24.255 210.355 24.685 211.140 ;
        RECT 24.705 210.415 26.075 211.225 ;
        RECT 26.085 210.415 31.595 211.225 ;
        RECT 31.605 210.415 37.115 211.225 ;
        RECT 37.135 210.355 37.565 211.140 ;
        RECT 37.585 210.415 38.955 211.225 ;
        RECT 38.965 210.415 44.475 211.225 ;
        RECT 44.485 210.415 49.995 211.225 ;
        RECT 50.015 210.355 50.445 211.140 ;
        RECT 50.465 210.415 51.835 211.225 ;
        RECT 51.845 210.415 57.355 211.225 ;
        RECT 57.365 210.415 62.875 211.225 ;
        RECT 62.895 210.355 63.325 211.140 ;
        RECT 63.345 210.415 64.715 211.225 ;
        RECT 64.725 210.415 70.235 211.225 ;
        RECT 70.245 210.415 75.755 211.225 ;
        RECT 75.775 210.355 76.205 211.140 ;
        RECT 76.225 210.415 77.595 211.225 ;
        RECT 77.605 210.415 83.115 211.225 ;
        RECT 83.125 210.415 88.635 211.225 ;
        RECT 88.655 210.355 89.085 211.140 ;
        RECT 89.105 210.415 90.475 211.225 ;
        RECT 90.485 210.415 95.995 211.225 ;
        RECT 96.005 210.415 101.515 211.225 ;
        RECT 101.535 210.355 101.965 211.140 ;
        RECT 101.985 210.415 103.355 211.225 ;
        RECT 103.365 210.415 108.875 211.225 ;
        RECT 108.885 210.415 114.395 211.225 ;
        RECT 114.415 210.355 114.845 211.140 ;
        RECT 115.325 210.415 120.835 211.225 ;
        RECT 120.845 210.415 126.355 211.225 ;
        RECT 126.365 210.415 127.735 211.225 ;
      LAYER nwell ;
        RECT 14.390 207.195 127.930 210.025 ;
      LAYER pwell ;
        RECT 14.585 205.995 15.955 206.805 ;
        RECT 15.965 205.995 18.715 206.805 ;
        RECT 18.725 205.995 24.235 206.805 ;
        RECT 24.255 206.080 24.685 206.865 ;
        RECT 25.165 205.995 27.915 206.805 ;
        RECT 27.925 205.995 33.435 206.805 ;
        RECT 33.445 205.995 38.955 206.805 ;
        RECT 38.965 205.995 44.475 206.805 ;
        RECT 44.485 205.995 49.995 206.805 ;
        RECT 50.015 206.080 50.445 206.865 ;
        RECT 50.465 205.995 55.975 206.805 ;
        RECT 55.985 205.995 61.495 206.805 ;
        RECT 61.505 205.995 67.015 206.805 ;
        RECT 67.025 205.995 72.535 206.805 ;
        RECT 72.555 205.995 73.905 206.905 ;
        RECT 74.410 206.675 75.755 206.905 ;
        RECT 73.925 205.995 75.755 206.675 ;
        RECT 75.775 206.080 76.205 206.865 ;
        RECT 77.145 205.995 80.255 206.905 ;
        RECT 81.285 205.995 84.955 206.805 ;
        RECT 84.965 205.995 90.475 206.805 ;
        RECT 90.485 205.995 95.995 206.805 ;
        RECT 96.005 205.995 101.515 206.805 ;
        RECT 101.535 206.080 101.965 206.865 ;
        RECT 102.445 205.995 104.275 206.805 ;
        RECT 104.285 205.995 109.795 206.805 ;
        RECT 109.805 205.995 115.315 206.805 ;
        RECT 115.325 205.995 120.835 206.805 ;
        RECT 120.845 205.995 126.355 206.805 ;
        RECT 126.365 205.995 127.735 206.805 ;
        RECT 14.725 205.785 14.895 205.995 ;
        RECT 16.565 205.830 16.725 205.940 ;
        RECT 18.405 205.805 18.575 205.995 ;
        RECT 20.245 205.785 20.415 205.975 ;
        RECT 23.925 205.805 24.095 205.995 ;
        RECT 24.900 205.835 25.020 205.945 ;
        RECT 25.765 205.785 25.935 205.975 ;
        RECT 27.605 205.805 27.775 205.995 ;
        RECT 31.285 205.785 31.455 205.975 ;
        RECT 33.125 205.805 33.295 205.995 ;
        RECT 36.805 205.785 36.975 205.975 ;
        RECT 37.780 205.835 37.900 205.945 ;
        RECT 38.645 205.805 38.815 205.995 ;
        RECT 40.485 205.785 40.655 205.975 ;
        RECT 44.165 205.805 44.335 205.995 ;
        RECT 46.005 205.785 46.175 205.975 ;
        RECT 49.685 205.805 49.855 205.995 ;
        RECT 51.525 205.785 51.695 205.975 ;
        RECT 55.665 205.805 55.835 205.995 ;
        RECT 57.045 205.785 57.215 205.975 ;
        RECT 61.185 205.805 61.355 205.995 ;
        RECT 62.565 205.785 62.735 205.975 ;
        RECT 64.405 205.785 64.575 205.975 ;
        RECT 65.785 205.785 65.955 205.975 ;
        RECT 66.705 205.805 66.875 205.995 ;
        RECT 67.165 205.785 67.335 205.975 ;
        RECT 72.225 205.805 72.395 205.995 ;
        RECT 72.685 205.805 72.855 205.995 ;
        RECT 74.065 205.805 74.235 205.995 ;
        RECT 76.825 205.840 76.985 205.950 ;
        RECT 77.285 205.785 77.455 205.975 ;
        RECT 80.045 205.805 80.215 205.995 ;
        RECT 80.965 205.840 81.125 205.950 ;
        RECT 84.645 205.805 84.815 205.995 ;
        RECT 86.485 205.785 86.655 205.975 ;
        RECT 88.325 205.785 88.495 205.975 ;
        RECT 89.300 205.835 89.420 205.945 ;
        RECT 90.165 205.805 90.335 205.995 ;
        RECT 92.005 205.785 92.175 205.975 ;
        RECT 95.685 205.805 95.855 205.995 ;
        RECT 97.525 205.785 97.695 205.975 ;
        RECT 101.205 205.805 101.375 205.995 ;
        RECT 102.180 205.835 102.300 205.945 ;
        RECT 103.045 205.785 103.215 205.975 ;
        RECT 103.965 205.805 104.135 205.995 ;
        RECT 108.565 205.785 108.735 205.975 ;
        RECT 109.485 205.805 109.655 205.995 ;
        RECT 114.085 205.785 114.255 205.975 ;
        RECT 115.005 205.945 115.175 205.995 ;
        RECT 115.005 205.835 115.180 205.945 ;
        RECT 115.005 205.805 115.175 205.835 ;
        RECT 120.525 205.785 120.695 205.995 ;
        RECT 126.045 205.785 126.215 205.995 ;
        RECT 127.425 205.785 127.595 205.995 ;
        RECT 14.585 204.975 15.955 205.785 ;
        RECT 16.885 204.975 20.555 205.785 ;
        RECT 20.565 204.975 26.075 205.785 ;
        RECT 26.085 204.975 31.595 205.785 ;
        RECT 31.605 204.975 37.115 205.785 ;
        RECT 37.135 204.915 37.565 205.700 ;
        RECT 38.045 204.975 40.795 205.785 ;
        RECT 40.805 204.975 46.315 205.785 ;
        RECT 46.325 204.975 51.835 205.785 ;
        RECT 51.845 204.975 57.355 205.785 ;
        RECT 57.365 204.975 62.875 205.785 ;
        RECT 62.895 204.915 63.325 205.700 ;
        RECT 63.345 204.975 64.715 205.785 ;
        RECT 64.735 204.875 66.085 205.785 ;
        RECT 67.035 204.875 68.385 205.785 ;
        RECT 68.405 205.105 77.595 205.785 ;
        RECT 77.605 205.105 86.795 205.785 ;
        RECT 68.405 204.875 69.325 205.105 ;
        RECT 72.155 204.885 73.085 205.105 ;
        RECT 77.605 204.875 78.525 205.105 ;
        RECT 81.355 204.885 82.285 205.105 ;
        RECT 86.805 204.975 88.635 205.785 ;
        RECT 88.655 204.915 89.085 205.700 ;
        RECT 89.565 204.975 92.315 205.785 ;
        RECT 92.325 204.975 97.835 205.785 ;
        RECT 97.845 204.975 103.355 205.785 ;
        RECT 103.365 204.975 108.875 205.785 ;
        RECT 108.885 204.975 114.395 205.785 ;
        RECT 114.415 204.915 114.845 205.700 ;
        RECT 115.325 204.975 120.835 205.785 ;
        RECT 120.845 204.975 126.355 205.785 ;
        RECT 126.365 204.975 127.735 205.785 ;
      LAYER nwell ;
        RECT 14.390 201.755 127.930 204.585 ;
      LAYER pwell ;
        RECT 14.585 200.555 15.955 201.365 ;
        RECT 15.965 200.555 18.715 201.365 ;
        RECT 18.725 200.555 24.235 201.365 ;
        RECT 24.255 200.640 24.685 201.425 ;
        RECT 25.165 200.555 27.915 201.365 ;
        RECT 27.925 200.555 33.435 201.365 ;
        RECT 33.445 200.555 38.955 201.365 ;
        RECT 38.965 200.555 44.475 201.365 ;
        RECT 44.485 200.555 49.995 201.365 ;
        RECT 50.015 200.640 50.445 201.425 ;
        RECT 50.465 200.555 54.135 201.365 ;
        RECT 54.145 200.555 59.655 201.365 ;
        RECT 64.175 201.235 65.105 201.455 ;
        RECT 67.825 201.235 70.035 201.465 ;
        RECT 59.665 200.555 70.035 201.235 ;
        RECT 70.245 201.235 71.175 201.465 ;
        RECT 70.245 200.555 73.915 201.235 ;
        RECT 73.925 200.555 75.755 201.235 ;
        RECT 75.775 200.640 76.205 201.425 ;
        RECT 76.685 201.235 77.605 201.465 ;
        RECT 79.445 201.235 80.365 201.465 ;
        RECT 83.195 201.235 84.125 201.455 ;
        RECT 76.685 200.555 78.975 201.235 ;
        RECT 79.445 200.555 88.635 201.235 ;
        RECT 88.645 200.555 90.475 201.365 ;
        RECT 90.485 200.555 95.995 201.365 ;
        RECT 96.005 200.555 101.515 201.365 ;
        RECT 101.535 200.640 101.965 201.425 ;
        RECT 102.445 200.555 104.275 201.365 ;
        RECT 104.285 200.555 109.795 201.365 ;
        RECT 109.805 200.555 115.315 201.365 ;
        RECT 115.325 200.555 120.835 201.365 ;
        RECT 120.845 200.555 126.355 201.365 ;
        RECT 126.365 200.555 127.735 201.365 ;
        RECT 14.725 200.345 14.895 200.555 ;
        RECT 16.565 200.390 16.725 200.500 ;
        RECT 18.405 200.365 18.575 200.555 ;
        RECT 20.245 200.345 20.415 200.535 ;
        RECT 23.925 200.365 24.095 200.555 ;
        RECT 24.900 200.395 25.020 200.505 ;
        RECT 25.765 200.345 25.935 200.535 ;
        RECT 27.605 200.365 27.775 200.555 ;
        RECT 31.285 200.345 31.455 200.535 ;
        RECT 33.125 200.365 33.295 200.555 ;
        RECT 36.805 200.345 36.975 200.535 ;
        RECT 37.780 200.395 37.900 200.505 ;
        RECT 38.645 200.365 38.815 200.555 ;
        RECT 40.485 200.345 40.655 200.535 ;
        RECT 44.165 200.365 44.335 200.555 ;
        RECT 46.005 200.345 46.175 200.535 ;
        RECT 49.685 200.365 49.855 200.555 ;
        RECT 51.525 200.345 51.695 200.535 ;
        RECT 53.825 200.365 53.995 200.555 ;
        RECT 57.045 200.345 57.215 200.535 ;
        RECT 59.345 200.365 59.515 200.555 ;
        RECT 59.805 200.365 59.975 200.555 ;
        RECT 62.565 200.345 62.735 200.535 ;
        RECT 63.540 200.395 63.660 200.505 ;
        RECT 67.165 200.345 67.335 200.535 ;
        RECT 68.545 200.345 68.715 200.535 ;
        RECT 70.385 200.345 70.555 200.535 ;
        RECT 73.605 200.365 73.775 200.555 ;
        RECT 74.985 200.345 75.155 200.535 ;
        RECT 75.445 200.365 75.615 200.555 ;
        RECT 76.420 200.395 76.540 200.505 ;
        RECT 78.665 200.345 78.835 200.555 ;
        RECT 79.180 200.395 79.300 200.505 ;
        RECT 80.965 200.365 81.135 200.535 ;
        RECT 80.965 200.345 81.130 200.365 ;
        RECT 82.350 200.345 82.520 200.535 ;
        RECT 82.805 200.345 82.975 200.535 ;
        RECT 84.185 200.345 84.355 200.535 ;
        RECT 86.485 200.345 86.655 200.535 ;
        RECT 88.325 200.345 88.495 200.555 ;
        RECT 89.300 200.395 89.420 200.505 ;
        RECT 90.165 200.365 90.335 200.555 ;
        RECT 91.085 200.345 91.255 200.535 ;
        RECT 95.685 200.365 95.855 200.555 ;
        RECT 96.605 200.345 96.775 200.535 ;
        RECT 101.205 200.365 101.375 200.555 ;
        RECT 102.180 200.395 102.300 200.505 ;
        RECT 103.965 200.365 104.135 200.555 ;
        RECT 105.805 200.345 105.975 200.535 ;
        RECT 108.565 200.345 108.735 200.535 ;
        RECT 109.485 200.365 109.655 200.555 ;
        RECT 114.085 200.345 114.255 200.535 ;
        RECT 115.005 200.505 115.175 200.555 ;
        RECT 115.005 200.395 115.180 200.505 ;
        RECT 115.005 200.365 115.175 200.395 ;
        RECT 120.525 200.345 120.695 200.555 ;
        RECT 126.045 200.345 126.215 200.555 ;
        RECT 127.425 200.345 127.595 200.555 ;
        RECT 14.585 199.535 15.955 200.345 ;
        RECT 16.885 199.535 20.555 200.345 ;
        RECT 20.565 199.535 26.075 200.345 ;
        RECT 26.085 199.535 31.595 200.345 ;
        RECT 31.605 199.535 37.115 200.345 ;
        RECT 37.135 199.475 37.565 200.260 ;
        RECT 38.045 199.535 40.795 200.345 ;
        RECT 40.805 199.535 46.315 200.345 ;
        RECT 46.325 199.535 51.835 200.345 ;
        RECT 51.845 199.535 57.355 200.345 ;
        RECT 57.365 199.535 62.875 200.345 ;
        RECT 62.895 199.475 63.325 200.260 ;
        RECT 63.805 199.535 67.475 200.345 ;
        RECT 67.485 199.565 68.855 200.345 ;
        RECT 68.865 199.665 70.695 200.345 ;
        RECT 70.715 200.305 71.635 200.345 ;
        RECT 70.705 200.115 71.635 200.305 ;
        RECT 73.725 200.115 75.295 200.345 ;
        RECT 70.705 199.755 75.295 200.115 ;
        RECT 70.715 199.665 75.295 199.755 ;
        RECT 75.400 199.665 78.865 200.345 ;
        RECT 79.295 199.665 81.130 200.345 ;
        RECT 70.715 199.435 73.715 199.665 ;
        RECT 75.400 199.435 76.320 199.665 ;
        RECT 79.295 199.435 80.225 199.665 ;
        RECT 81.285 199.435 82.635 200.345 ;
        RECT 82.665 199.565 84.035 200.345 ;
        RECT 84.055 199.435 85.405 200.345 ;
        RECT 85.435 199.435 86.785 200.345 ;
        RECT 86.805 199.535 88.635 200.345 ;
        RECT 88.655 199.475 89.085 200.260 ;
        RECT 89.565 199.535 91.395 200.345 ;
        RECT 91.405 199.535 96.915 200.345 ;
        RECT 96.925 199.665 106.115 200.345 ;
        RECT 96.925 199.435 97.845 199.665 ;
        RECT 100.675 199.445 101.605 199.665 ;
        RECT 106.125 199.535 108.875 200.345 ;
        RECT 108.885 199.535 114.395 200.345 ;
        RECT 114.415 199.475 114.845 200.260 ;
        RECT 115.325 199.535 120.835 200.345 ;
        RECT 120.845 199.535 126.355 200.345 ;
        RECT 126.365 199.535 127.735 200.345 ;
      LAYER nwell ;
        RECT 14.390 196.315 127.930 199.145 ;
      LAYER pwell ;
        RECT 14.585 195.115 15.955 195.925 ;
        RECT 15.965 195.115 18.715 195.925 ;
        RECT 18.725 195.115 24.235 195.925 ;
        RECT 24.255 195.200 24.685 195.985 ;
        RECT 25.165 195.115 27.915 195.925 ;
        RECT 27.925 195.115 33.435 195.925 ;
        RECT 33.445 195.115 38.955 195.925 ;
        RECT 38.965 195.115 44.475 195.925 ;
        RECT 44.485 195.115 49.995 195.925 ;
        RECT 50.015 195.200 50.445 195.985 ;
        RECT 50.925 195.115 52.755 195.925 ;
        RECT 52.775 195.115 54.125 196.025 ;
        RECT 56.800 195.795 57.720 196.025 ;
        RECT 54.255 195.115 57.720 195.795 ;
        RECT 57.825 195.115 63.335 195.925 ;
        RECT 63.345 195.115 68.855 195.925 ;
        RECT 68.865 195.795 69.785 196.025 ;
        RECT 68.865 195.115 71.155 195.795 ;
        RECT 71.165 195.115 74.085 196.025 ;
        RECT 74.385 195.115 75.755 195.925 ;
        RECT 75.775 195.200 76.205 195.985 ;
        RECT 76.225 195.115 79.895 195.925 ;
        RECT 79.905 195.115 85.415 195.925 ;
        RECT 85.795 195.915 86.715 196.025 ;
        RECT 85.795 195.795 88.130 195.915 ;
        RECT 92.795 195.795 93.715 196.015 ;
        RECT 85.795 195.115 95.075 195.795 ;
        RECT 95.085 195.115 97.835 195.925 ;
        RECT 100.500 195.795 101.420 196.025 ;
        RECT 97.955 195.115 101.420 195.795 ;
        RECT 101.535 195.200 101.965 195.985 ;
        RECT 101.985 195.115 104.735 195.925 ;
        RECT 104.745 195.115 110.255 195.925 ;
        RECT 110.265 195.795 111.185 196.025 ;
        RECT 114.015 195.795 114.945 196.015 ;
        RECT 110.265 195.115 119.455 195.795 ;
        RECT 119.465 195.115 120.835 195.925 ;
        RECT 120.845 195.115 126.355 195.925 ;
        RECT 126.365 195.115 127.735 195.925 ;
        RECT 14.725 194.905 14.895 195.115 ;
        RECT 16.565 194.950 16.725 195.060 ;
        RECT 18.405 194.925 18.575 195.115 ;
        RECT 20.245 194.905 20.415 195.095 ;
        RECT 23.925 194.925 24.095 195.115 ;
        RECT 24.900 194.955 25.020 195.065 ;
        RECT 25.765 194.905 25.935 195.095 ;
        RECT 27.605 194.925 27.775 195.115 ;
        RECT 31.285 194.905 31.455 195.095 ;
        RECT 33.125 194.925 33.295 195.115 ;
        RECT 36.805 194.905 36.975 195.095 ;
        RECT 38.185 194.950 38.345 195.060 ;
        RECT 38.645 194.925 38.815 195.115 ;
        RECT 41.865 194.905 42.035 195.095 ;
        RECT 44.165 194.925 44.335 195.115 ;
        RECT 47.385 194.905 47.555 195.095 ;
        RECT 48.765 194.905 48.935 195.095 ;
        RECT 49.225 194.905 49.395 195.095 ;
        RECT 49.685 194.925 49.855 195.115 ;
        RECT 50.660 194.955 50.780 195.065 ;
        RECT 52.445 194.925 52.615 195.115 ;
        RECT 53.825 194.925 53.995 195.115 ;
        RECT 54.285 194.925 54.455 195.115 ;
        RECT 58.885 194.950 59.045 195.060 ;
        RECT 62.565 194.905 62.735 195.095 ;
        RECT 63.025 194.925 63.195 195.115 ;
        RECT 64.865 194.905 65.035 195.095 ;
        RECT 66.245 194.905 66.415 195.095 ;
        RECT 66.760 194.955 66.880 195.065 ;
        RECT 68.545 194.905 68.715 195.115 ;
        RECT 14.585 194.095 15.955 194.905 ;
        RECT 16.885 194.095 20.555 194.905 ;
        RECT 20.565 194.095 26.075 194.905 ;
        RECT 26.085 194.095 31.595 194.905 ;
        RECT 31.605 194.095 37.115 194.905 ;
        RECT 37.135 194.035 37.565 194.820 ;
        RECT 38.505 194.095 42.175 194.905 ;
        RECT 42.185 194.095 47.695 194.905 ;
        RECT 47.715 193.995 49.065 194.905 ;
        RECT 49.085 194.225 58.275 194.905 ;
        RECT 53.595 194.005 54.525 194.225 ;
        RECT 57.355 193.995 58.275 194.225 ;
        RECT 59.205 194.095 62.875 194.905 ;
        RECT 62.895 194.035 63.325 194.820 ;
        RECT 63.345 194.095 65.175 194.905 ;
        RECT 65.195 193.995 66.545 194.905 ;
        RECT 67.025 194.095 68.855 194.905 ;
        RECT 69.005 194.875 69.175 195.095 ;
        RECT 70.845 194.925 71.015 195.115 ;
        RECT 71.310 194.925 71.480 195.115 ;
        RECT 71.130 194.875 72.075 194.905 ;
        RECT 69.005 194.675 72.075 194.875 ;
        RECT 68.865 194.195 72.075 194.675 ;
        RECT 68.865 193.995 69.795 194.195 ;
        RECT 71.130 193.995 72.075 194.195 ;
        RECT 72.085 194.875 73.030 194.905 ;
        RECT 74.985 194.875 75.155 195.095 ;
        RECT 75.445 194.925 75.615 195.115 ;
        RECT 78.665 194.905 78.835 195.095 ;
        RECT 79.585 194.925 79.755 195.115 ;
        RECT 84.185 194.905 84.355 195.095 ;
        RECT 85.105 194.925 85.275 195.115 ;
        RECT 88.050 194.905 88.220 195.095 ;
        RECT 90.165 194.905 90.335 195.095 ;
        RECT 92.925 194.905 93.095 195.095 ;
        RECT 93.385 194.905 93.555 195.095 ;
        RECT 94.765 194.905 94.935 195.115 ;
        RECT 97.525 194.925 97.695 195.115 ;
        RECT 97.985 194.925 98.155 195.115 ;
        RECT 104.425 194.925 104.595 195.115 ;
        RECT 104.885 194.905 105.055 195.095 ;
        RECT 108.565 194.905 108.735 195.095 ;
        RECT 109.025 194.905 109.195 195.095 ;
        RECT 109.945 194.925 110.115 195.115 ;
        RECT 113.810 194.905 113.980 195.095 ;
        RECT 115.925 194.905 116.095 195.095 ;
        RECT 116.845 194.950 117.005 195.060 ;
        RECT 119.145 194.925 119.315 195.115 ;
        RECT 120.525 194.905 120.695 195.115 ;
        RECT 126.045 194.905 126.215 195.115 ;
        RECT 127.425 194.905 127.595 195.115 ;
        RECT 72.085 194.675 75.155 194.875 ;
        RECT 72.085 194.195 75.295 194.675 ;
        RECT 72.085 193.995 73.030 194.195 ;
        RECT 74.365 193.995 75.295 194.195 ;
        RECT 75.305 194.095 78.975 194.905 ;
        RECT 78.985 194.095 84.495 194.905 ;
        RECT 84.735 194.225 88.635 194.905 ;
        RECT 87.705 193.995 88.635 194.225 ;
        RECT 88.655 194.035 89.085 194.820 ;
        RECT 89.115 193.995 90.465 194.905 ;
        RECT 90.485 194.095 93.235 194.905 ;
        RECT 93.255 193.995 94.605 194.905 ;
        RECT 94.625 194.225 103.730 194.905 ;
        RECT 103.825 194.095 105.195 194.905 ;
        RECT 105.205 194.095 108.875 194.905 ;
        RECT 108.895 193.995 110.245 194.905 ;
        RECT 110.495 194.225 114.395 194.905 ;
        RECT 113.465 193.995 114.395 194.225 ;
        RECT 114.415 194.035 114.845 194.820 ;
        RECT 114.875 193.995 116.225 194.905 ;
        RECT 117.165 194.095 120.835 194.905 ;
        RECT 120.845 194.095 126.355 194.905 ;
        RECT 126.365 194.095 127.735 194.905 ;
      LAYER nwell ;
        RECT 14.390 190.875 127.930 193.705 ;
      LAYER pwell ;
        RECT 14.585 189.675 15.955 190.485 ;
        RECT 15.965 189.675 18.715 190.485 ;
        RECT 18.725 189.675 24.235 190.485 ;
        RECT 24.255 189.760 24.685 190.545 ;
        RECT 25.165 189.675 30.675 190.485 ;
        RECT 30.685 189.675 36.195 190.485 ;
        RECT 36.575 190.475 37.495 190.585 ;
        RECT 36.575 190.355 38.910 190.475 ;
        RECT 43.575 190.355 44.495 190.575 ;
        RECT 49.065 190.355 49.995 190.585 ;
        RECT 36.575 189.675 45.855 190.355 ;
        RECT 46.095 189.675 49.995 190.355 ;
        RECT 50.015 189.760 50.445 190.545 ;
        RECT 50.925 189.675 52.295 190.455 ;
        RECT 52.305 190.355 53.225 190.585 ;
        RECT 56.055 190.355 56.985 190.575 ;
        RECT 61.545 190.355 62.885 190.585 ;
        RECT 65.715 190.355 66.645 190.575 ;
        RECT 52.305 189.675 61.495 190.355 ;
        RECT 61.545 189.675 71.155 190.355 ;
        RECT 71.165 189.675 74.275 190.585 ;
        RECT 74.385 189.675 75.755 190.485 ;
        RECT 75.775 189.760 76.205 190.545 ;
        RECT 76.225 189.675 78.515 190.585 ;
        RECT 79.445 189.675 83.115 190.485 ;
        RECT 83.495 190.475 84.415 190.585 ;
        RECT 83.495 190.355 85.830 190.475 ;
        RECT 90.495 190.355 91.415 190.575 ;
        RECT 83.495 189.675 92.775 190.355 ;
        RECT 92.785 189.675 94.155 190.455 ;
        RECT 100.585 190.355 101.515 190.585 ;
        RECT 94.545 189.675 96.970 190.355 ;
        RECT 97.615 189.675 101.515 190.355 ;
        RECT 101.535 189.760 101.965 190.545 ;
        RECT 101.985 189.675 103.355 190.455 ;
        RECT 103.365 189.675 104.735 190.485 ;
        RECT 107.945 190.355 108.875 190.585 ;
        RECT 104.975 189.675 108.875 190.355 ;
        RECT 108.885 190.355 109.805 190.585 ;
        RECT 112.635 190.355 113.565 190.575 ;
        RECT 108.885 189.675 118.075 190.355 ;
        RECT 118.085 189.675 119.455 190.455 ;
        RECT 119.465 189.675 120.835 190.485 ;
        RECT 120.845 189.675 126.355 190.485 ;
        RECT 126.365 189.675 127.735 190.485 ;
        RECT 14.725 189.465 14.895 189.675 ;
        RECT 16.160 189.515 16.280 189.625 ;
        RECT 17.945 189.465 18.115 189.655 ;
        RECT 18.405 189.485 18.575 189.675 ;
        RECT 23.465 189.465 23.635 189.655 ;
        RECT 23.925 189.485 24.095 189.675 ;
        RECT 24.900 189.515 25.020 189.625 ;
        RECT 28.985 189.465 29.155 189.655 ;
        RECT 30.365 189.465 30.535 189.675 ;
        RECT 31.745 189.465 31.915 189.655 ;
        RECT 35.425 189.465 35.595 189.655 ;
        RECT 35.885 189.465 36.055 189.675 ;
        RECT 45.545 189.485 45.715 189.675 ;
        RECT 46.465 189.465 46.635 189.655 ;
        RECT 49.410 189.485 49.580 189.675 ;
        RECT 50.660 189.515 50.780 189.625 ;
        RECT 51.985 189.485 52.155 189.675 ;
        RECT 55.665 189.465 55.835 189.655 ;
        RECT 59.530 189.465 59.700 189.655 ;
        RECT 61.185 189.465 61.355 189.675 ;
        RECT 62.565 189.465 62.735 189.655 ;
        RECT 63.540 189.515 63.660 189.625 ;
        RECT 63.945 189.465 64.115 189.655 ;
        RECT 69.925 189.465 70.095 189.655 ;
        RECT 70.845 189.485 71.015 189.675 ;
        RECT 74.065 189.485 74.235 189.675 ;
        RECT 75.445 189.465 75.615 189.675 ;
        RECT 76.370 189.485 76.540 189.675 ;
        RECT 79.125 189.520 79.285 189.630 ;
        RECT 80.965 189.465 81.135 189.655 ;
        RECT 82.805 189.485 82.975 189.675 ;
        RECT 86.485 189.465 86.655 189.655 ;
        RECT 87.865 189.465 88.035 189.655 ;
        RECT 88.380 189.515 88.500 189.625 ;
        RECT 89.245 189.465 89.415 189.655 ;
        RECT 92.005 189.465 92.175 189.655 ;
        RECT 92.465 189.485 92.635 189.675 ;
        RECT 92.925 189.485 93.095 189.675 ;
        RECT 97.065 189.485 97.235 189.655 ;
        RECT 97.525 189.465 97.695 189.655 ;
        RECT 100.930 189.485 101.100 189.675 ;
        RECT 102.125 189.485 102.295 189.675 ;
        RECT 104.425 189.485 104.595 189.675 ;
        RECT 106.725 189.465 106.895 189.655 ;
        RECT 108.290 189.485 108.460 189.675 ;
        RECT 110.405 189.465 110.575 189.655 ;
        RECT 110.920 189.515 111.040 189.625 ;
        RECT 112.705 189.465 112.875 189.655 ;
        RECT 113.165 189.465 113.335 189.655 ;
        RECT 115.060 189.515 115.180 189.625 ;
        RECT 117.765 189.485 117.935 189.675 ;
        RECT 119.145 189.485 119.315 189.675 ;
        RECT 120.525 189.465 120.695 189.675 ;
        RECT 126.045 189.465 126.215 189.675 ;
        RECT 127.425 189.465 127.595 189.675 ;
        RECT 14.585 188.655 15.955 189.465 ;
        RECT 16.425 188.655 18.255 189.465 ;
        RECT 18.265 188.655 23.775 189.465 ;
        RECT 23.785 188.655 29.295 189.465 ;
        RECT 29.315 188.555 30.665 189.465 ;
        RECT 30.685 188.655 32.055 189.465 ;
        RECT 32.065 188.655 35.735 189.465 ;
        RECT 35.755 188.555 37.105 189.465 ;
        RECT 37.135 188.595 37.565 189.380 ;
        RECT 37.585 188.785 46.775 189.465 ;
        RECT 46.870 188.785 55.975 189.465 ;
        RECT 56.215 188.785 60.115 189.465 ;
        RECT 37.585 188.555 38.505 188.785 ;
        RECT 41.335 188.565 42.265 188.785 ;
        RECT 59.185 188.555 60.115 188.785 ;
        RECT 60.125 188.685 61.495 189.465 ;
        RECT 61.505 188.655 62.875 189.465 ;
        RECT 62.895 188.595 63.325 189.380 ;
        RECT 63.915 188.785 67.380 189.465 ;
        RECT 66.460 188.555 67.380 188.785 ;
        RECT 67.485 188.655 70.235 189.465 ;
        RECT 70.245 188.655 75.755 189.465 ;
        RECT 75.765 188.655 81.275 189.465 ;
        RECT 81.285 188.655 86.795 189.465 ;
        RECT 86.815 188.555 88.165 189.465 ;
        RECT 88.655 188.595 89.085 189.380 ;
        RECT 89.105 188.685 90.475 189.465 ;
        RECT 90.485 188.655 92.315 189.465 ;
        RECT 92.325 188.655 97.835 189.465 ;
        RECT 97.845 188.785 107.035 189.465 ;
        RECT 107.140 188.785 110.605 189.465 ;
        RECT 97.845 188.555 98.765 188.785 ;
        RECT 101.595 188.565 102.525 188.785 ;
        RECT 107.140 188.555 108.060 188.785 ;
        RECT 111.185 188.655 113.015 189.465 ;
        RECT 113.025 188.685 114.395 189.465 ;
        RECT 114.415 188.595 114.845 189.380 ;
        RECT 115.325 188.655 120.835 189.465 ;
        RECT 120.845 188.655 126.355 189.465 ;
        RECT 126.365 188.655 127.735 189.465 ;
      LAYER nwell ;
        RECT 14.390 185.435 127.930 188.265 ;
      LAYER pwell ;
        RECT 14.585 184.235 15.955 185.045 ;
        RECT 15.965 184.235 18.715 185.045 ;
        RECT 18.725 184.235 24.235 185.045 ;
        RECT 24.255 184.320 24.685 185.105 ;
        RECT 24.705 184.235 26.075 185.045 ;
        RECT 26.085 184.915 27.005 185.145 ;
        RECT 29.835 184.915 30.765 185.135 ;
        RECT 26.085 184.235 35.275 184.915 ;
        RECT 35.745 184.235 38.495 185.045 ;
        RECT 38.515 184.235 39.865 185.145 ;
        RECT 43.085 184.915 44.015 185.145 ;
        RECT 40.115 184.235 44.015 184.915 ;
        RECT 44.025 184.915 44.955 185.145 ;
        RECT 44.025 184.235 47.925 184.915 ;
        RECT 48.635 184.235 49.985 185.145 ;
        RECT 50.015 184.320 50.445 185.105 ;
        RECT 50.465 184.915 51.385 185.145 ;
        RECT 54.215 184.915 55.145 185.135 ;
        RECT 50.465 184.235 59.655 184.915 ;
        RECT 60.125 184.235 65.635 185.045 ;
        RECT 65.645 184.235 71.155 185.045 ;
        RECT 71.175 184.915 74.175 185.145 ;
        RECT 71.175 184.825 75.755 184.915 ;
        RECT 71.165 184.465 75.755 184.825 ;
        RECT 71.165 184.275 72.095 184.465 ;
        RECT 71.175 184.235 72.095 184.275 ;
        RECT 74.185 184.235 75.755 184.465 ;
        RECT 75.775 184.320 76.205 185.105 ;
        RECT 76.225 184.235 78.975 185.045 ;
        RECT 78.985 184.235 84.495 185.045 ;
        RECT 87.705 184.915 88.635 185.145 ;
        RECT 84.735 184.235 88.635 184.915 ;
        RECT 88.645 184.235 94.155 185.045 ;
        RECT 96.820 184.915 97.740 185.145 ;
        RECT 94.275 184.235 97.740 184.915 ;
        RECT 98.765 184.235 100.135 185.015 ;
        RECT 100.155 184.235 101.505 185.145 ;
        RECT 101.535 184.320 101.965 185.105 ;
        RECT 102.540 184.915 103.460 185.145 ;
        RECT 109.240 184.915 110.160 185.145 ;
        RECT 112.920 184.915 113.840 185.145 ;
        RECT 102.540 184.235 106.005 184.915 ;
        RECT 106.695 184.235 110.160 184.915 ;
        RECT 110.375 184.235 113.840 184.915 ;
        RECT 113.945 184.235 115.315 185.045 ;
        RECT 115.325 184.235 120.835 185.045 ;
        RECT 120.845 184.235 126.355 185.045 ;
        RECT 126.365 184.235 127.735 185.045 ;
        RECT 14.725 184.025 14.895 184.235 ;
        RECT 16.160 184.075 16.280 184.185 ;
        RECT 18.405 184.045 18.575 184.235 ;
        RECT 21.625 184.025 21.795 184.215 ;
        RECT 22.085 184.025 22.255 184.215 ;
        RECT 23.925 184.045 24.095 184.235 ;
        RECT 25.765 184.045 25.935 184.235 ;
        RECT 26.685 184.025 26.855 184.215 ;
        RECT 27.145 184.025 27.315 184.215 ;
        RECT 31.100 184.025 31.270 184.215 ;
        RECT 34.965 184.185 35.135 184.235 ;
        RECT 34.965 184.075 35.140 184.185 ;
        RECT 35.480 184.075 35.600 184.185 ;
        RECT 34.965 184.045 35.135 184.075 ;
        RECT 36.805 184.025 36.975 184.215 ;
        RECT 37.725 184.025 37.895 184.215 ;
        RECT 38.185 184.045 38.355 184.235 ;
        RECT 38.645 184.045 38.815 184.235 ;
        RECT 41.405 184.025 41.575 184.215 ;
        RECT 43.430 184.045 43.600 184.235 ;
        RECT 44.440 184.045 44.610 184.235 ;
        RECT 45.085 184.025 45.255 184.215 ;
        RECT 48.360 184.075 48.480 184.185 ;
        RECT 48.765 184.045 48.935 184.235 ;
        RECT 49.685 184.025 49.855 184.215 ;
        RECT 51.065 184.025 51.235 184.215 ;
        RECT 51.525 184.025 51.695 184.215 ;
        RECT 55.665 184.025 55.835 184.215 ;
        RECT 56.180 184.075 56.300 184.185 ;
        RECT 58.885 184.025 59.055 184.215 ;
        RECT 59.345 184.045 59.515 184.235 ;
        RECT 59.860 184.075 59.980 184.185 ;
        RECT 60.265 184.025 60.435 184.215 ;
        RECT 60.780 184.075 60.900 184.185 ;
        RECT 62.565 184.025 62.735 184.215 ;
        RECT 63.540 184.075 63.660 184.185 ;
        RECT 65.325 184.045 65.495 184.235 ;
        RECT 66.245 184.025 66.415 184.215 ;
        RECT 66.705 184.045 66.875 184.215 ;
        RECT 66.805 184.025 66.875 184.045 ;
        RECT 69.925 184.025 70.095 184.215 ;
        RECT 70.845 184.045 71.015 184.235 ;
        RECT 75.445 184.045 75.615 184.235 ;
        RECT 78.205 184.045 78.375 184.215 ;
        RECT 78.665 184.045 78.835 184.235 ;
        RECT 79.125 184.070 79.285 184.180 ;
        RECT 84.185 184.045 84.355 184.235 ;
        RECT 88.050 184.045 88.220 184.235 ;
        RECT 78.205 184.025 78.275 184.045 ;
        RECT 88.325 184.025 88.495 184.215 ;
        RECT 90.165 184.025 90.335 184.215 ;
        RECT 91.545 184.025 91.715 184.215 ;
        RECT 93.845 184.045 94.015 184.235 ;
        RECT 94.305 184.045 94.475 184.235 ;
        RECT 95.225 184.025 95.395 184.215 ;
        RECT 98.445 184.080 98.605 184.190 ;
        RECT 98.905 184.045 99.075 184.235 ;
        RECT 99.090 184.025 99.260 184.215 ;
        RECT 100.285 184.045 100.455 184.235 ;
        RECT 102.125 184.185 102.295 184.215 ;
        RECT 102.125 184.075 102.300 184.185 ;
        RECT 102.125 184.025 102.295 184.075 ;
        RECT 105.805 184.045 105.975 184.235 ;
        RECT 106.725 184.215 106.895 184.235 ;
        RECT 105.990 184.025 106.160 184.215 ;
        RECT 106.320 184.075 106.440 184.185 ;
        RECT 106.725 184.045 106.900 184.215 ;
        RECT 110.405 184.045 110.575 184.235 ;
        RECT 106.730 184.025 106.900 184.045 ;
        RECT 113.810 184.025 113.980 184.215 ;
        RECT 115.005 184.045 115.175 184.235 ;
        RECT 115.465 184.070 115.625 184.180 ;
        RECT 120.525 184.045 120.695 184.235 ;
        RECT 124.665 184.025 124.835 184.215 ;
        RECT 126.045 184.025 126.215 184.235 ;
        RECT 127.425 184.025 127.595 184.235 ;
        RECT 14.585 183.215 15.955 184.025 ;
        RECT 16.425 183.215 21.935 184.025 ;
        RECT 21.945 183.245 23.315 184.025 ;
        RECT 23.420 183.345 26.885 184.025 ;
        RECT 27.115 183.345 30.580 184.025 ;
        RECT 23.420 183.115 24.340 183.345 ;
        RECT 29.660 183.115 30.580 183.345 ;
        RECT 30.685 183.345 34.585 184.025 ;
        RECT 30.685 183.115 31.615 183.345 ;
        RECT 35.285 183.215 37.115 184.025 ;
        RECT 37.135 183.155 37.565 183.940 ;
        RECT 37.695 183.345 41.160 184.025 ;
        RECT 41.375 183.345 44.840 184.025 ;
        RECT 45.055 183.345 48.520 184.025 ;
        RECT 40.240 183.115 41.160 183.345 ;
        RECT 43.920 183.115 44.840 183.345 ;
        RECT 47.600 183.115 48.520 183.345 ;
        RECT 48.625 183.245 49.995 184.025 ;
        RECT 50.005 183.245 51.375 184.025 ;
        RECT 51.385 183.245 52.755 184.025 ;
        RECT 52.765 183.115 55.925 184.025 ;
        RECT 56.445 183.215 59.195 184.025 ;
        RECT 59.215 183.115 60.565 184.025 ;
        RECT 61.045 183.215 62.875 184.025 ;
        RECT 62.895 183.155 63.325 183.940 ;
        RECT 63.805 183.215 66.555 184.025 ;
        RECT 66.805 183.795 69.075 184.025 ;
        RECT 69.785 183.795 74.210 184.025 ;
        RECT 76.005 183.795 78.275 184.025 ;
        RECT 66.805 183.115 69.560 183.795 ;
        RECT 69.785 183.115 75.150 183.795 ;
        RECT 75.520 183.115 78.275 183.795 ;
        RECT 79.445 183.345 88.635 184.025 ;
        RECT 79.445 183.115 80.365 183.345 ;
        RECT 83.195 183.125 84.125 183.345 ;
        RECT 88.655 183.155 89.085 183.940 ;
        RECT 89.115 183.115 90.465 184.025 ;
        RECT 90.485 183.215 91.855 184.025 ;
        RECT 91.865 183.215 95.535 184.025 ;
        RECT 95.775 183.345 99.675 184.025 ;
        RECT 98.745 183.115 99.675 183.345 ;
        RECT 99.685 183.215 102.435 184.025 ;
        RECT 102.675 183.345 106.575 184.025 ;
        RECT 105.645 183.115 106.575 183.345 ;
        RECT 106.585 183.115 110.060 184.025 ;
        RECT 110.495 183.345 114.395 184.025 ;
        RECT 113.465 183.115 114.395 183.345 ;
        RECT 114.415 183.155 114.845 183.940 ;
        RECT 115.785 183.345 124.975 184.025 ;
        RECT 115.785 183.115 116.705 183.345 ;
        RECT 119.535 183.125 120.465 183.345 ;
        RECT 124.985 183.215 126.355 184.025 ;
        RECT 126.365 183.215 127.735 184.025 ;
      LAYER nwell ;
        RECT 14.390 179.995 127.930 182.825 ;
      LAYER pwell ;
        RECT 14.585 178.795 15.955 179.605 ;
        RECT 15.965 178.795 18.715 179.605 ;
        RECT 18.725 178.795 24.235 179.605 ;
        RECT 24.255 178.880 24.685 179.665 ;
        RECT 29.215 179.475 30.145 179.695 ;
        RECT 32.975 179.475 33.895 179.705 ;
        RECT 24.705 178.795 33.895 179.475 ;
        RECT 34.000 179.475 34.920 179.705 ;
        RECT 34.000 178.795 37.465 179.475 ;
        RECT 38.045 178.795 41.520 179.705 ;
        RECT 42.185 178.795 45.660 179.705 ;
        RECT 49.065 179.475 49.995 179.705 ;
        RECT 46.095 178.795 49.995 179.475 ;
        RECT 50.015 178.880 50.445 179.665 ;
        RECT 53.120 179.475 54.040 179.705 ;
        RECT 50.575 178.795 54.040 179.475 ;
        RECT 54.145 178.795 55.975 179.605 ;
        RECT 55.985 179.475 56.915 179.705 ;
        RECT 55.985 178.795 59.885 179.475 ;
        RECT 60.135 178.795 62.875 179.475 ;
        RECT 62.885 178.795 65.635 179.605 ;
        RECT 65.655 178.795 67.005 179.705 ;
        RECT 67.025 179.475 68.370 179.705 ;
        RECT 67.025 178.795 68.855 179.475 ;
        RECT 68.865 178.795 71.605 179.475 ;
        RECT 71.865 179.025 74.620 179.705 ;
        RECT 71.865 178.795 74.135 179.025 ;
        RECT 75.775 178.880 76.205 179.665 ;
        RECT 78.880 179.475 79.800 179.705 ;
        RECT 76.335 178.795 79.800 179.475 ;
        RECT 80.100 178.795 83.575 179.705 ;
        RECT 83.585 178.795 85.415 179.605 ;
        RECT 88.625 179.475 89.555 179.705 ;
        RECT 85.655 178.795 89.555 179.475 ;
        RECT 89.565 178.795 90.935 179.575 ;
        RECT 90.955 178.795 92.305 179.705 ;
        RECT 92.325 179.475 93.245 179.705 ;
        RECT 96.075 179.475 97.005 179.695 ;
        RECT 92.325 178.795 101.515 179.475 ;
        RECT 101.535 178.880 101.965 179.665 ;
        RECT 102.080 179.475 103.000 179.705 ;
        RECT 105.760 179.475 106.680 179.705 ;
        RECT 102.080 178.795 105.545 179.475 ;
        RECT 105.760 178.795 109.225 179.475 ;
        RECT 109.815 178.795 111.165 179.705 ;
        RECT 111.185 179.475 112.105 179.705 ;
        RECT 114.935 179.475 115.865 179.695 ;
        RECT 111.185 178.795 120.375 179.475 ;
        RECT 120.395 178.795 121.745 179.705 ;
        RECT 121.765 178.795 123.135 179.575 ;
        RECT 123.605 178.795 126.355 179.605 ;
        RECT 126.365 178.795 127.735 179.605 ;
        RECT 14.725 178.585 14.895 178.795 ;
        RECT 18.405 178.605 18.575 178.795 ;
        RECT 19.325 178.585 19.495 178.775 ;
        RECT 23.925 178.605 24.095 178.795 ;
        RECT 24.845 178.585 25.015 178.795 ;
        RECT 26.225 178.585 26.395 178.775 ;
        RECT 26.685 178.585 26.855 178.775 ;
        RECT 36.805 178.585 36.975 178.775 ;
        RECT 37.265 178.605 37.435 178.795 ;
        RECT 37.780 178.635 37.900 178.745 ;
        RECT 38.190 178.605 38.360 178.795 ;
        RECT 41.130 178.585 41.300 178.775 ;
        RECT 41.920 178.635 42.040 178.745 ;
        RECT 42.330 178.740 42.500 178.795 ;
        RECT 42.325 178.630 42.500 178.740 ;
        RECT 42.330 178.605 42.500 178.630 ;
        RECT 42.785 178.585 42.955 178.775 ;
        RECT 49.410 178.605 49.580 178.795 ;
        RECT 49.680 178.585 49.850 178.775 ;
        RECT 50.145 178.585 50.315 178.775 ;
        RECT 50.605 178.605 50.775 178.795 ;
        RECT 55.665 178.605 55.835 178.795 ;
        RECT 56.400 178.605 56.570 178.795 ;
        RECT 62.565 178.585 62.735 178.795 ;
        RECT 64.405 178.585 64.575 178.775 ;
        RECT 65.325 178.605 65.495 178.795 ;
        RECT 65.785 178.605 65.955 178.795 ;
        RECT 67.165 178.585 67.335 178.775 ;
        RECT 68.545 178.605 68.715 178.795 ;
        RECT 69.005 178.585 69.175 178.795 ;
        RECT 71.865 178.775 71.935 178.795 ;
        RECT 69.465 178.585 69.635 178.775 ;
        RECT 71.305 178.585 71.475 178.775 ;
        RECT 71.765 178.605 71.935 178.775 ;
        RECT 75.445 178.585 75.615 178.775 ;
        RECT 75.960 178.635 76.080 178.745 ;
        RECT 76.365 178.605 76.535 178.795 ;
        RECT 79.580 178.585 79.750 178.775 ;
        RECT 80.050 178.585 80.220 178.775 ;
        RECT 83.260 178.605 83.430 178.795 ;
        RECT 84.645 178.585 84.815 178.775 ;
        RECT 85.105 178.585 85.275 178.795 ;
        RECT 88.970 178.605 89.140 178.795 ;
        RECT 90.625 178.605 90.795 178.795 ;
        RECT 91.085 178.605 91.255 178.795 ;
        RECT 92.465 178.585 92.635 178.775 ;
        RECT 97.985 178.585 98.155 178.775 ;
        RECT 101.205 178.605 101.375 178.795 ;
        RECT 101.660 178.585 101.830 178.775 ;
        RECT 103.045 178.585 103.215 178.775 ;
        RECT 104.425 178.585 104.595 178.775 ;
        RECT 104.890 178.585 105.060 178.775 ;
        RECT 105.345 178.605 105.515 178.795 ;
        RECT 109.025 178.605 109.195 178.795 ;
        RECT 109.540 178.635 109.660 178.745 ;
        RECT 109.945 178.585 110.115 178.795 ;
        RECT 113.810 178.585 113.980 178.775 ;
        RECT 116.385 178.585 116.555 178.775 ;
        RECT 116.845 178.585 117.015 178.775 ;
        RECT 120.065 178.605 120.235 178.795 ;
        RECT 120.525 178.585 120.695 178.795 ;
        RECT 121.905 178.605 122.075 178.795 ;
        RECT 123.340 178.635 123.460 178.745 ;
        RECT 126.045 178.585 126.215 178.795 ;
        RECT 127.425 178.585 127.595 178.795 ;
        RECT 14.585 177.775 15.955 178.585 ;
        RECT 15.965 177.775 19.635 178.585 ;
        RECT 19.645 177.775 25.155 178.585 ;
        RECT 25.175 177.675 26.525 178.585 ;
        RECT 26.555 177.675 27.905 178.585 ;
        RECT 27.925 177.905 37.115 178.585 ;
        RECT 27.925 177.675 28.845 177.905 ;
        RECT 31.675 177.685 32.605 177.905 ;
        RECT 37.135 177.715 37.565 178.500 ;
        RECT 37.815 177.905 41.715 178.585 ;
        RECT 42.755 177.905 46.220 178.585 ;
        RECT 40.785 177.675 41.715 177.905 ;
        RECT 45.300 177.675 46.220 177.905 ;
        RECT 46.520 177.675 49.995 178.585 ;
        RECT 50.115 177.905 53.580 178.585 ;
        RECT 52.660 177.675 53.580 177.905 ;
        RECT 53.685 177.905 62.875 178.585 ;
        RECT 53.685 177.675 54.605 177.905 ;
        RECT 57.435 177.685 58.365 177.905 ;
        RECT 62.895 177.715 63.325 178.500 ;
        RECT 63.345 177.805 64.715 178.585 ;
        RECT 64.725 177.775 67.475 178.585 ;
        RECT 67.485 177.905 69.315 178.585 ;
        RECT 69.325 177.905 71.155 178.585 ;
        RECT 71.165 177.905 72.995 178.585 ;
        RECT 67.485 177.675 68.830 177.905 ;
        RECT 69.810 177.675 71.155 177.905 ;
        RECT 71.650 177.675 72.995 177.905 ;
        RECT 73.035 177.675 75.755 178.585 ;
        RECT 76.420 177.675 79.895 178.585 ;
        RECT 79.905 177.675 83.380 178.585 ;
        RECT 83.585 177.775 84.955 178.585 ;
        RECT 85.075 177.905 88.540 178.585 ;
        RECT 87.620 177.675 88.540 177.905 ;
        RECT 88.655 177.715 89.085 178.500 ;
        RECT 89.105 177.775 92.775 178.585 ;
        RECT 92.785 177.775 98.295 178.585 ;
        RECT 98.500 177.675 101.975 178.585 ;
        RECT 101.985 177.805 103.355 178.585 ;
        RECT 103.365 177.775 104.735 178.585 ;
        RECT 104.745 177.675 108.220 178.585 ;
        RECT 108.425 177.775 110.255 178.585 ;
        RECT 110.495 177.905 114.395 178.585 ;
        RECT 113.465 177.675 114.395 177.905 ;
        RECT 114.415 177.715 114.845 178.500 ;
        RECT 114.865 177.775 116.695 178.585 ;
        RECT 116.705 177.805 118.075 178.585 ;
        RECT 118.085 177.775 120.835 178.585 ;
        RECT 120.845 177.775 126.355 178.585 ;
        RECT 126.365 177.775 127.735 178.585 ;
      LAYER nwell ;
        RECT 14.390 174.555 127.930 177.385 ;
      LAYER pwell ;
        RECT 14.585 173.355 15.955 174.165 ;
        RECT 15.965 173.355 18.715 174.165 ;
        RECT 18.725 173.355 24.235 174.165 ;
        RECT 24.255 173.440 24.685 174.225 ;
        RECT 25.625 173.355 26.995 174.135 ;
        RECT 29.660 174.035 30.580 174.265 ;
        RECT 27.115 173.355 30.580 174.035 ;
        RECT 30.685 174.035 31.615 174.265 ;
        RECT 30.685 173.355 34.585 174.035 ;
        RECT 35.480 173.355 38.955 174.265 ;
        RECT 38.965 173.355 42.440 174.265 ;
        RECT 42.840 173.355 46.315 174.265 ;
        RECT 48.980 174.035 49.900 174.265 ;
        RECT 46.435 173.355 49.900 174.035 ;
        RECT 50.015 173.440 50.445 174.225 ;
        RECT 50.465 173.355 53.215 174.165 ;
        RECT 56.425 174.035 57.355 174.265 ;
        RECT 53.455 173.355 57.355 174.035 ;
        RECT 57.365 174.035 58.285 174.265 ;
        RECT 61.115 174.035 62.045 174.255 ;
        RECT 57.365 173.355 66.555 174.035 ;
        RECT 66.565 173.355 68.395 174.165 ;
        RECT 68.405 173.355 71.015 174.265 ;
        RECT 71.165 174.035 72.510 174.265 ;
        RECT 71.165 173.355 72.995 174.035 ;
        RECT 73.005 173.355 75.755 174.165 ;
        RECT 75.775 173.440 76.205 174.225 ;
        RECT 77.145 173.355 80.815 174.165 ;
        RECT 80.825 173.355 84.300 174.265 ;
        RECT 84.965 173.355 90.475 174.165 ;
        RECT 90.485 173.355 95.995 174.165 ;
        RECT 96.005 173.355 101.515 174.165 ;
        RECT 101.535 173.440 101.965 174.225 ;
        RECT 101.985 173.355 103.815 174.165 ;
        RECT 104.020 173.355 107.495 174.265 ;
        RECT 107.505 173.355 110.980 174.265 ;
        RECT 111.185 173.355 112.555 174.165 ;
        RECT 112.565 173.355 118.075 174.165 ;
        RECT 118.095 173.355 119.445 174.265 ;
        RECT 119.465 173.355 120.835 174.165 ;
        RECT 120.845 173.355 126.355 174.165 ;
        RECT 126.365 173.355 127.735 174.165 ;
        RECT 14.725 173.145 14.895 173.355 ;
        RECT 16.565 173.190 16.725 173.300 ;
        RECT 18.405 173.165 18.575 173.355 ;
        RECT 20.245 173.145 20.415 173.335 ;
        RECT 23.925 173.165 24.095 173.355 ;
        RECT 25.305 173.200 25.465 173.310 ;
        RECT 25.765 173.145 25.935 173.335 ;
        RECT 26.685 173.165 26.855 173.355 ;
        RECT 27.145 173.165 27.315 173.355 ;
        RECT 31.100 173.165 31.270 173.355 ;
        RECT 31.285 173.145 31.455 173.335 ;
        RECT 35.020 173.195 35.140 173.305 ;
        RECT 36.805 173.145 36.975 173.335 ;
        RECT 37.730 173.145 37.900 173.335 ;
        RECT 38.640 173.165 38.810 173.355 ;
        RECT 39.110 173.165 39.280 173.355 ;
        RECT 41.460 173.195 41.580 173.305 ;
        RECT 42.785 173.145 42.955 173.335 ;
        RECT 43.705 173.190 43.865 173.300 ;
        RECT 44.170 173.145 44.340 173.335 ;
        RECT 46.000 173.165 46.170 173.355 ;
        RECT 46.465 173.165 46.635 173.355 ;
        RECT 47.850 173.145 48.020 173.335 ;
        RECT 51.530 173.145 51.700 173.335 ;
        RECT 52.905 173.165 53.075 173.355 ;
        RECT 56.125 173.145 56.295 173.335 ;
        RECT 56.770 173.165 56.940 173.355 ;
        RECT 59.805 173.145 59.975 173.335 ;
        RECT 61.185 173.145 61.355 173.335 ;
        RECT 61.645 173.145 61.815 173.335 ;
        RECT 63.540 173.195 63.660 173.305 ;
        RECT 65.325 173.145 65.495 173.335 ;
        RECT 66.245 173.165 66.415 173.355 ;
        RECT 68.085 173.165 68.255 173.355 ;
        RECT 68.550 173.165 68.720 173.355 ;
        RECT 70.845 173.145 71.015 173.335 ;
        RECT 72.685 173.165 72.855 173.355 ;
        RECT 75.445 173.165 75.615 173.355 ;
        RECT 76.365 173.145 76.535 173.335 ;
        RECT 76.825 173.200 76.985 173.310 ;
        RECT 80.505 173.165 80.675 173.355 ;
        RECT 80.970 173.165 81.140 173.355 ;
        RECT 81.885 173.145 82.055 173.335 ;
        RECT 82.350 173.145 82.520 173.335 ;
        RECT 84.700 173.195 84.820 173.305 ;
        RECT 85.105 173.145 85.275 173.335 ;
        RECT 89.300 173.195 89.420 173.305 ;
        RECT 89.705 173.145 89.875 173.335 ;
        RECT 90.165 173.165 90.335 173.355 ;
        RECT 95.685 173.165 95.855 173.355 ;
        RECT 99.825 173.145 99.995 173.335 ;
        RECT 100.745 173.190 100.905 173.300 ;
        RECT 101.205 173.165 101.375 173.355 ;
        RECT 103.505 173.165 103.675 173.355 ;
        RECT 106.265 173.145 106.435 173.335 ;
        RECT 107.180 173.165 107.350 173.355 ;
        RECT 107.650 173.335 107.820 173.355 ;
        RECT 107.645 173.165 107.820 173.335 ;
        RECT 107.645 173.145 107.815 173.165 ;
        RECT 111.320 173.145 111.490 173.335 ;
        RECT 112.245 173.165 112.415 173.355 ;
        RECT 112.705 173.145 112.875 173.335 ;
        RECT 113.165 173.145 113.335 173.335 ;
        RECT 115.465 173.190 115.625 173.300 ;
        RECT 117.765 173.165 117.935 173.355 ;
        RECT 118.225 173.165 118.395 173.355 ;
        RECT 120.525 173.165 120.695 173.355 ;
        RECT 124.665 173.145 124.835 173.335 ;
        RECT 126.045 173.145 126.215 173.355 ;
        RECT 127.425 173.145 127.595 173.355 ;
        RECT 14.585 172.335 15.955 173.145 ;
        RECT 16.885 172.335 20.555 173.145 ;
        RECT 20.565 172.335 26.075 173.145 ;
        RECT 26.085 172.335 31.595 173.145 ;
        RECT 31.605 172.335 37.115 173.145 ;
        RECT 37.135 172.275 37.565 173.060 ;
        RECT 37.585 172.235 41.060 173.145 ;
        RECT 41.725 172.365 43.095 173.145 ;
        RECT 44.025 172.235 47.500 173.145 ;
        RECT 47.705 172.235 51.180 173.145 ;
        RECT 51.385 172.235 54.860 173.145 ;
        RECT 55.065 172.335 56.435 173.145 ;
        RECT 56.445 172.335 60.115 173.145 ;
        RECT 60.135 172.235 61.485 173.145 ;
        RECT 61.505 172.365 62.875 173.145 ;
        RECT 62.895 172.275 63.325 173.060 ;
        RECT 63.805 172.335 65.635 173.145 ;
        RECT 65.645 172.335 71.155 173.145 ;
        RECT 71.165 172.335 76.675 173.145 ;
        RECT 76.685 172.335 82.195 173.145 ;
        RECT 82.205 172.235 84.815 173.145 ;
        RECT 85.075 172.465 88.540 173.145 ;
        RECT 87.620 172.235 88.540 172.465 ;
        RECT 88.655 172.275 89.085 173.060 ;
        RECT 89.575 172.235 90.925 173.145 ;
        RECT 90.945 172.465 100.135 173.145 ;
        RECT 90.945 172.235 91.865 172.465 ;
        RECT 94.695 172.245 95.625 172.465 ;
        RECT 101.065 172.335 106.575 173.145 ;
        RECT 106.595 172.235 107.945 173.145 ;
        RECT 108.160 172.235 111.635 173.145 ;
        RECT 111.645 172.335 113.015 173.145 ;
        RECT 113.035 172.235 114.385 173.145 ;
        RECT 114.415 172.275 114.845 173.060 ;
        RECT 115.785 172.465 124.975 173.145 ;
        RECT 115.785 172.235 116.705 172.465 ;
        RECT 119.535 172.245 120.465 172.465 ;
        RECT 124.985 172.335 126.355 173.145 ;
        RECT 126.365 172.335 127.735 173.145 ;
      LAYER nwell ;
        RECT 14.390 169.115 127.930 171.945 ;
      LAYER pwell ;
        RECT 14.585 167.915 15.955 168.725 ;
        RECT 15.965 167.915 18.715 168.725 ;
        RECT 18.725 167.915 24.235 168.725 ;
        RECT 24.255 168.000 24.685 168.785 ;
        RECT 25.165 167.915 26.995 168.725 ;
        RECT 27.015 167.915 28.365 168.825 ;
        RECT 28.845 167.915 32.515 168.725 ;
        RECT 32.535 167.915 33.885 168.825 ;
        RECT 33.905 167.915 35.275 168.725 ;
        RECT 35.370 167.915 44.475 168.595 ;
        RECT 44.485 167.915 49.995 168.725 ;
        RECT 50.015 168.000 50.445 168.785 ;
        RECT 50.465 167.915 51.835 168.725 ;
        RECT 51.845 167.915 57.355 168.725 ;
        RECT 57.365 167.915 62.875 168.725 ;
        RECT 62.885 167.915 68.395 168.725 ;
        RECT 68.405 168.595 69.750 168.825 ;
        RECT 70.245 168.595 71.590 168.825 ;
        RECT 68.405 167.915 70.235 168.595 ;
        RECT 70.245 167.915 72.075 168.595 ;
        RECT 72.085 167.915 75.755 168.725 ;
        RECT 75.775 168.000 76.205 168.785 ;
        RECT 79.425 168.595 80.355 168.825 ;
        RECT 76.455 167.915 80.355 168.595 ;
        RECT 80.735 168.715 81.655 168.825 ;
        RECT 80.735 168.595 83.070 168.715 ;
        RECT 87.735 168.595 88.655 168.815 ;
        RECT 80.735 167.915 90.015 168.595 ;
        RECT 90.025 167.915 91.395 168.725 ;
        RECT 94.605 168.595 95.535 168.825 ;
        RECT 91.635 167.915 95.535 168.595 ;
        RECT 96.005 167.915 97.375 168.695 ;
        RECT 97.845 167.915 101.515 168.725 ;
        RECT 101.535 168.000 101.965 168.785 ;
        RECT 102.905 168.595 103.825 168.825 ;
        RECT 106.655 168.595 107.585 168.815 ;
        RECT 112.565 168.595 113.495 168.825 ;
        RECT 116.800 168.595 117.720 168.825 ;
        RECT 102.905 167.915 112.095 168.595 ;
        RECT 112.565 167.915 116.465 168.595 ;
        RECT 116.800 167.915 120.265 168.595 ;
        RECT 120.385 167.915 121.755 168.695 ;
        RECT 121.765 167.915 123.595 168.595 ;
        RECT 123.605 167.915 126.355 168.725 ;
        RECT 126.365 167.915 127.735 168.725 ;
        RECT 14.725 167.705 14.895 167.915 ;
        RECT 17.485 167.705 17.655 167.895 ;
        RECT 18.405 167.725 18.575 167.915 ;
        RECT 23.005 167.705 23.175 167.895 ;
        RECT 23.465 167.705 23.635 167.895 ;
        RECT 23.925 167.725 24.095 167.915 ;
        RECT 24.900 167.755 25.020 167.865 ;
        RECT 26.685 167.725 26.855 167.915 ;
        RECT 27.145 167.725 27.315 167.915 ;
        RECT 28.580 167.755 28.700 167.865 ;
        RECT 32.205 167.725 32.375 167.915 ;
        RECT 33.585 167.705 33.755 167.915 ;
        RECT 34.965 167.725 35.135 167.915 ;
        RECT 36.805 167.705 36.975 167.895 ;
        RECT 37.725 167.705 37.895 167.895 ;
        RECT 39.105 167.705 39.275 167.895 ;
        RECT 44.165 167.725 44.335 167.915 ;
        RECT 46.005 167.705 46.175 167.895 ;
        RECT 46.925 167.750 47.085 167.860 ;
        RECT 49.685 167.725 49.855 167.915 ;
        RECT 51.525 167.725 51.695 167.915 ;
        RECT 56.125 167.705 56.295 167.895 ;
        RECT 57.045 167.725 57.215 167.915 ;
        RECT 62.565 167.895 62.735 167.915 ;
        RECT 57.965 167.705 58.135 167.895 ;
        RECT 59.345 167.705 59.515 167.895 ;
        RECT 59.860 167.755 59.980 167.865 ;
        RECT 62.560 167.725 62.735 167.895 ;
        RECT 62.560 167.705 62.730 167.725 ;
        RECT 64.865 167.705 65.035 167.895 ;
        RECT 67.625 167.705 67.795 167.895 ;
        RECT 68.085 167.705 68.255 167.915 ;
        RECT 69.925 167.725 70.095 167.915 ;
        RECT 70.845 167.705 71.015 167.895 ;
        RECT 71.765 167.725 71.935 167.915 ;
        RECT 74.985 167.705 75.155 167.895 ;
        RECT 75.445 167.725 75.615 167.915 ;
        RECT 79.770 167.725 79.940 167.915 ;
        RECT 84.645 167.705 84.815 167.895 ;
        RECT 86.025 167.705 86.195 167.895 ;
        RECT 87.405 167.705 87.575 167.895 ;
        RECT 88.325 167.750 88.485 167.860 ;
        RECT 89.300 167.755 89.420 167.865 ;
        RECT 89.705 167.725 89.875 167.915 ;
        RECT 91.085 167.725 91.255 167.915 ;
        RECT 92.925 167.705 93.095 167.895 ;
        RECT 94.950 167.725 95.120 167.915 ;
        RECT 95.740 167.755 95.860 167.865 ;
        RECT 96.145 167.725 96.315 167.915 ;
        RECT 96.790 167.705 96.960 167.895 ;
        RECT 97.580 167.755 97.700 167.865 ;
        RECT 101.205 167.725 101.375 167.915 ;
        RECT 102.585 167.760 102.745 167.870 ;
        RECT 106.725 167.705 106.895 167.895 ;
        RECT 107.185 167.705 107.355 167.895 ;
        RECT 110.865 167.705 111.035 167.895 ;
        RECT 111.785 167.725 111.955 167.915 ;
        RECT 112.300 167.755 112.420 167.865 ;
        RECT 112.980 167.725 113.150 167.915 ;
        RECT 115.465 167.750 115.625 167.860 ;
        RECT 120.065 167.725 120.235 167.915 ;
        RECT 120.525 167.725 120.695 167.915 ;
        RECT 123.285 167.725 123.455 167.915 ;
        RECT 124.665 167.705 124.835 167.895 ;
        RECT 126.045 167.705 126.215 167.915 ;
        RECT 127.425 167.705 127.595 167.915 ;
        RECT 14.585 166.895 15.955 167.705 ;
        RECT 15.965 166.895 17.795 167.705 ;
        RECT 17.805 166.895 23.315 167.705 ;
        RECT 23.325 167.025 32.515 167.705 ;
        RECT 27.835 166.805 28.765 167.025 ;
        RECT 31.595 166.795 32.515 167.025 ;
        RECT 32.525 166.925 33.895 167.705 ;
        RECT 33.905 166.795 37.065 167.705 ;
        RECT 37.135 166.835 37.565 167.620 ;
        RECT 37.595 166.795 38.945 167.705 ;
        RECT 39.075 167.025 42.540 167.705 ;
        RECT 41.620 166.795 42.540 167.025 ;
        RECT 42.740 167.025 46.205 167.705 ;
        RECT 47.245 167.025 56.435 167.705 ;
        RECT 42.740 166.795 43.660 167.025 ;
        RECT 47.245 166.795 48.165 167.025 ;
        RECT 50.995 166.805 51.925 167.025 ;
        RECT 56.445 166.895 58.275 167.705 ;
        RECT 58.295 166.795 59.645 167.705 ;
        RECT 60.265 166.795 62.875 167.705 ;
        RECT 62.895 166.835 63.325 167.620 ;
        RECT 63.345 166.895 65.175 167.705 ;
        RECT 65.195 167.025 67.935 167.705 ;
        RECT 67.945 167.025 70.685 167.705 ;
        RECT 70.705 166.795 73.425 167.705 ;
        RECT 73.465 166.895 75.295 167.705 ;
        RECT 75.675 167.025 84.955 167.705 ;
        RECT 75.675 166.905 78.010 167.025 ;
        RECT 75.675 166.795 76.595 166.905 ;
        RECT 82.675 166.805 83.595 167.025 ;
        RECT 84.975 166.795 86.325 167.705 ;
        RECT 86.355 166.795 87.705 167.705 ;
        RECT 88.655 166.835 89.085 167.620 ;
        RECT 89.565 166.895 93.235 167.705 ;
        RECT 93.475 167.025 97.375 167.705 ;
        RECT 96.445 166.795 97.375 167.025 ;
        RECT 97.755 167.025 107.035 167.705 ;
        RECT 107.155 167.025 110.620 167.705 ;
        RECT 110.835 167.025 114.300 167.705 ;
        RECT 97.755 166.905 100.090 167.025 ;
        RECT 97.755 166.795 98.675 166.905 ;
        RECT 104.755 166.805 105.675 167.025 ;
        RECT 109.700 166.795 110.620 167.025 ;
        RECT 113.380 166.795 114.300 167.025 ;
        RECT 114.415 166.835 114.845 167.620 ;
        RECT 115.785 167.025 124.975 167.705 ;
        RECT 115.785 166.795 116.705 167.025 ;
        RECT 119.535 166.805 120.465 167.025 ;
        RECT 124.985 166.895 126.355 167.705 ;
        RECT 126.365 166.895 127.735 167.705 ;
      LAYER nwell ;
        RECT 14.390 163.675 127.930 166.505 ;
      LAYER pwell ;
        RECT 14.585 162.475 15.955 163.285 ;
        RECT 15.965 162.475 18.715 163.285 ;
        RECT 18.725 162.475 24.235 163.285 ;
        RECT 24.255 162.560 24.685 163.345 ;
        RECT 25.625 162.475 26.995 163.255 ;
        RECT 31.515 163.155 32.445 163.375 ;
        RECT 35.275 163.155 36.195 163.385 ;
        RECT 27.005 162.475 36.195 163.155 ;
        RECT 36.205 163.155 37.125 163.385 ;
        RECT 39.955 163.155 40.885 163.375 ;
        RECT 48.980 163.155 49.900 163.385 ;
        RECT 36.205 162.475 45.395 163.155 ;
        RECT 46.435 162.475 49.900 163.155 ;
        RECT 50.015 162.560 50.445 163.345 ;
        RECT 50.475 162.475 51.825 163.385 ;
        RECT 51.845 162.475 53.675 163.285 ;
        RECT 53.685 162.475 55.055 163.255 ;
        RECT 55.065 163.155 55.985 163.385 ;
        RECT 58.815 163.155 59.745 163.375 ;
        RECT 55.065 162.475 64.255 163.155 ;
        RECT 64.405 162.475 67.015 163.385 ;
        RECT 67.035 162.475 69.775 163.155 ;
        RECT 70.245 162.475 75.755 163.285 ;
        RECT 75.775 162.560 76.205 163.345 ;
        RECT 76.225 162.475 78.055 163.285 ;
        RECT 81.265 163.155 82.195 163.385 ;
        RECT 78.295 162.475 82.195 163.155 ;
        RECT 82.205 162.475 83.575 163.255 ;
        RECT 83.585 162.475 85.415 163.285 ;
        RECT 85.425 162.475 86.795 163.255 ;
        RECT 86.805 162.475 92.315 163.285 ;
        RECT 92.410 162.475 101.515 163.155 ;
        RECT 101.535 162.560 101.965 163.345 ;
        RECT 105.185 163.155 106.115 163.385 ;
        RECT 102.215 162.475 106.115 163.155 ;
        RECT 106.585 163.155 107.515 163.385 ;
        RECT 106.585 162.475 110.485 163.155 ;
        RECT 110.865 162.475 113.475 163.385 ;
        RECT 113.485 163.155 114.405 163.385 ;
        RECT 117.235 163.155 118.165 163.375 ;
        RECT 113.485 162.475 122.675 163.155 ;
        RECT 122.685 162.475 124.055 163.255 ;
        RECT 124.525 162.475 126.355 163.285 ;
        RECT 126.365 162.475 127.735 163.285 ;
        RECT 14.725 162.265 14.895 162.475 ;
        RECT 17.485 162.265 17.655 162.455 ;
        RECT 18.405 162.285 18.575 162.475 ;
        RECT 23.925 162.285 24.095 162.475 ;
        RECT 25.305 162.320 25.465 162.430 ;
        RECT 26.685 162.285 26.855 162.475 ;
        RECT 27.145 162.265 27.315 162.475 ;
        RECT 27.880 162.265 28.050 162.455 ;
        RECT 32.665 162.265 32.835 162.455 ;
        RECT 33.400 162.265 33.570 162.455 ;
        RECT 37.780 162.315 37.900 162.425 ;
        RECT 39.565 162.265 39.735 162.455 ;
        RECT 40.025 162.265 40.195 162.455 ;
        RECT 43.980 162.265 44.150 162.455 ;
        RECT 45.085 162.285 45.255 162.475 ;
        RECT 46.005 162.320 46.165 162.430 ;
        RECT 46.465 162.285 46.635 162.475 ;
        RECT 48.765 162.265 48.935 162.455 ;
        RECT 49.500 162.265 49.670 162.455 ;
        RECT 51.525 162.285 51.695 162.475 ;
        RECT 53.365 162.285 53.535 162.475 ;
        RECT 53.825 162.285 53.995 162.475 ;
        RECT 56.770 162.265 56.940 162.455 ;
        RECT 57.560 162.315 57.680 162.425 ;
        RECT 59.345 162.265 59.515 162.455 ;
        RECT 59.805 162.265 59.975 162.455 ;
        RECT 62.565 162.265 62.735 162.455 ;
        RECT 63.945 162.285 64.115 162.475 ;
        RECT 64.405 162.265 64.575 162.455 ;
        RECT 66.245 162.265 66.415 162.455 ;
        RECT 66.700 162.285 66.870 162.475 ;
        RECT 68.085 162.265 68.255 162.455 ;
        RECT 68.545 162.265 68.715 162.455 ;
        RECT 69.465 162.285 69.635 162.475 ;
        RECT 69.980 162.315 70.100 162.425 ;
        RECT 70.385 162.265 70.555 162.455 ;
        RECT 72.280 162.315 72.400 162.425 ;
        RECT 74.985 162.265 75.155 162.455 ;
        RECT 75.445 162.285 75.615 162.475 ;
        RECT 77.745 162.285 77.915 162.475 ;
        RECT 80.505 162.265 80.675 162.455 ;
        RECT 81.610 162.285 81.780 162.475 ;
        RECT 81.885 162.265 82.055 162.455 ;
        RECT 82.345 162.285 82.515 162.475 ;
        RECT 85.105 162.285 85.275 162.475 ;
        RECT 85.565 162.285 85.735 162.475 ;
        RECT 85.750 162.265 85.920 162.455 ;
        RECT 86.485 162.265 86.655 162.455 ;
        RECT 88.325 162.310 88.485 162.420 ;
        RECT 89.300 162.315 89.420 162.425 ;
        RECT 92.005 162.285 92.175 162.475 ;
        RECT 98.905 162.265 99.075 162.455 ;
        RECT 101.205 162.285 101.375 162.475 ;
        RECT 102.125 162.265 102.295 162.455 ;
        RECT 102.585 162.265 102.755 162.455 ;
        RECT 105.530 162.285 105.700 162.475 ;
        RECT 106.320 162.315 106.440 162.425 ;
        RECT 106.725 162.265 106.895 162.455 ;
        RECT 107.000 162.285 107.170 162.475 ;
        RECT 113.160 162.285 113.330 162.475 ;
        RECT 113.810 162.265 113.980 162.455 ;
        RECT 118.410 162.265 118.580 162.455 ;
        RECT 119.145 162.265 119.315 162.455 ;
        RECT 120.580 162.315 120.700 162.425 ;
        RECT 120.985 162.265 121.155 162.455 ;
        RECT 122.365 162.425 122.535 162.475 ;
        RECT 122.365 162.315 122.540 162.425 ;
        RECT 122.365 162.285 122.535 162.315 ;
        RECT 123.745 162.285 123.915 162.475 ;
        RECT 124.260 162.315 124.380 162.425 ;
        RECT 126.045 162.265 126.215 162.475 ;
        RECT 127.425 162.265 127.595 162.475 ;
        RECT 14.585 161.455 15.955 162.265 ;
        RECT 15.965 161.455 17.795 162.265 ;
        RECT 18.175 161.585 27.455 162.265 ;
        RECT 27.465 161.585 31.365 162.265 ;
        RECT 18.175 161.465 20.510 161.585 ;
        RECT 18.175 161.355 19.095 161.465 ;
        RECT 25.175 161.365 26.095 161.585 ;
        RECT 27.465 161.355 28.395 161.585 ;
        RECT 31.605 161.455 32.975 162.265 ;
        RECT 32.985 161.585 36.885 162.265 ;
        RECT 32.985 161.355 33.915 161.585 ;
        RECT 37.135 161.395 37.565 162.180 ;
        RECT 38.045 161.455 39.875 162.265 ;
        RECT 39.995 161.585 43.460 162.265 ;
        RECT 42.540 161.355 43.460 161.585 ;
        RECT 43.565 161.585 47.465 162.265 ;
        RECT 43.565 161.355 44.495 161.585 ;
        RECT 47.705 161.485 49.075 162.265 ;
        RECT 49.085 161.585 52.985 162.265 ;
        RECT 53.455 161.585 57.355 162.265 ;
        RECT 49.085 161.355 50.015 161.585 ;
        RECT 56.425 161.355 57.355 161.585 ;
        RECT 57.825 161.455 59.655 162.265 ;
        RECT 59.665 161.485 61.035 162.265 ;
        RECT 61.045 161.455 62.875 162.265 ;
        RECT 62.895 161.395 63.325 162.180 ;
        RECT 63.345 161.455 64.715 162.265 ;
        RECT 64.725 161.585 66.555 162.265 ;
        RECT 66.565 161.585 68.395 162.265 ;
        RECT 68.405 161.585 70.235 162.265 ;
        RECT 70.245 161.585 72.075 162.265 ;
        RECT 64.725 161.355 66.070 161.585 ;
        RECT 66.565 161.355 67.910 161.585 ;
        RECT 68.890 161.355 70.235 161.585 ;
        RECT 70.730 161.355 72.075 161.585 ;
        RECT 72.545 161.455 75.295 162.265 ;
        RECT 75.305 161.455 80.815 162.265 ;
        RECT 80.835 161.355 82.185 162.265 ;
        RECT 82.435 161.585 86.335 162.265 ;
        RECT 85.405 161.355 86.335 161.585 ;
        RECT 86.345 161.485 87.715 162.265 ;
        RECT 88.655 161.395 89.085 162.180 ;
        RECT 89.935 161.585 99.215 162.265 ;
        RECT 89.935 161.465 92.270 161.585 ;
        RECT 89.935 161.355 90.855 161.465 ;
        RECT 96.935 161.365 97.855 161.585 ;
        RECT 99.225 161.355 102.385 162.265 ;
        RECT 102.555 161.585 106.020 162.265 ;
        RECT 106.695 161.585 110.160 162.265 ;
        RECT 110.495 161.585 114.395 162.265 ;
        RECT 105.100 161.355 106.020 161.585 ;
        RECT 109.240 161.355 110.160 161.585 ;
        RECT 113.465 161.355 114.395 161.585 ;
        RECT 114.415 161.395 114.845 162.180 ;
        RECT 115.095 161.585 118.995 162.265 ;
        RECT 118.065 161.355 118.995 161.585 ;
        RECT 119.015 161.355 120.365 162.265 ;
        RECT 120.845 161.485 122.215 162.265 ;
        RECT 122.685 161.455 126.355 162.265 ;
        RECT 126.365 161.455 127.735 162.265 ;
      LAYER nwell ;
        RECT 14.390 158.235 127.930 161.065 ;
      LAYER pwell ;
        RECT 14.585 157.035 15.955 157.845 ;
        RECT 15.965 157.035 17.335 157.845 ;
        RECT 17.355 157.035 18.705 157.945 ;
        RECT 18.735 157.035 20.085 157.945 ;
        RECT 23.305 157.715 24.235 157.945 ;
        RECT 20.335 157.035 24.235 157.715 ;
        RECT 24.255 157.120 24.685 157.905 ;
        RECT 24.705 157.035 26.075 157.815 ;
        RECT 26.085 157.035 27.915 157.845 ;
        RECT 30.580 157.715 31.500 157.945 ;
        RECT 34.260 157.715 35.180 157.945 ;
        RECT 28.035 157.035 31.500 157.715 ;
        RECT 31.715 157.035 35.180 157.715 ;
        RECT 35.285 157.035 38.955 157.845 ;
        RECT 39.160 157.035 42.635 157.945 ;
        RECT 42.840 157.035 46.315 157.945 ;
        RECT 48.980 157.715 49.900 157.945 ;
        RECT 46.435 157.035 49.900 157.715 ;
        RECT 50.015 157.120 50.445 157.905 ;
        RECT 50.465 157.035 53.940 157.945 ;
        RECT 54.605 157.035 60.115 157.845 ;
        RECT 60.135 157.035 61.485 157.945 ;
        RECT 61.645 157.035 64.255 157.945 ;
        RECT 64.725 157.035 68.395 157.845 ;
        RECT 68.890 157.715 70.235 157.945 ;
        RECT 70.730 157.715 72.075 157.945 ;
        RECT 68.405 157.035 70.235 157.715 ;
        RECT 70.245 157.035 72.075 157.715 ;
        RECT 72.280 157.035 75.755 157.945 ;
        RECT 75.775 157.120 76.205 157.905 ;
        RECT 76.880 157.035 80.355 157.945 ;
        RECT 81.195 157.835 82.115 157.945 ;
        RECT 81.195 157.715 83.530 157.835 ;
        RECT 88.195 157.715 89.115 157.935 ;
        RECT 81.195 157.035 90.475 157.715 ;
        RECT 90.945 157.035 92.775 157.845 ;
        RECT 92.795 157.035 94.145 157.945 ;
        RECT 94.625 157.035 96.455 157.845 ;
        RECT 96.465 157.035 97.835 157.815 ;
        RECT 97.845 157.035 99.675 157.845 ;
        RECT 99.695 157.035 101.045 157.945 ;
        RECT 101.535 157.120 101.965 157.905 ;
        RECT 102.445 157.035 104.275 157.845 ;
        RECT 104.285 157.035 105.655 157.815 ;
        RECT 105.665 157.035 107.035 157.815 ;
        RECT 107.965 157.035 111.440 157.945 ;
        RECT 112.565 157.035 116.235 157.845 ;
        RECT 118.900 157.715 119.820 157.945 ;
        RECT 116.355 157.035 119.820 157.715 ;
        RECT 120.845 157.035 126.355 157.845 ;
        RECT 126.365 157.035 127.735 157.845 ;
        RECT 14.725 156.825 14.895 157.035 ;
        RECT 16.565 156.870 16.725 156.980 ;
        RECT 17.025 156.845 17.195 157.035 ;
        RECT 18.405 156.845 18.575 157.035 ;
        RECT 18.865 156.845 19.035 157.035 ;
        RECT 23.650 156.845 23.820 157.035 ;
        RECT 24.845 156.845 25.015 157.035 ;
        RECT 26.225 156.825 26.395 157.015 ;
        RECT 27.605 156.825 27.775 157.035 ;
        RECT 28.065 156.845 28.235 157.035 ;
        RECT 28.985 156.825 29.155 157.015 ;
        RECT 31.745 156.845 31.915 157.035 ;
        RECT 32.665 156.825 32.835 157.015 ;
        RECT 36.530 156.825 36.700 157.015 ;
        RECT 37.780 156.875 37.900 156.985 ;
        RECT 38.645 156.845 38.815 157.035 ;
        RECT 39.565 156.825 39.735 157.015 ;
        RECT 40.030 156.825 40.200 157.015 ;
        RECT 42.320 156.845 42.490 157.035 ;
        RECT 43.710 156.825 43.880 157.015 ;
        RECT 46.000 156.845 46.170 157.035 ;
        RECT 46.465 156.845 46.635 157.035 ;
        RECT 47.390 156.825 47.560 157.015 ;
        RECT 50.610 156.845 50.780 157.035 ;
        RECT 51.120 156.875 51.240 156.985 ;
        RECT 52.905 156.825 53.075 157.015 ;
        RECT 54.340 156.875 54.460 156.985 ;
        RECT 59.805 156.845 59.975 157.035 ;
        RECT 61.185 156.845 61.355 157.035 ;
        RECT 62.565 156.825 62.735 157.015 ;
        RECT 63.540 156.875 63.660 156.985 ;
        RECT 63.940 156.845 64.110 157.035 ;
        RECT 64.460 156.875 64.580 156.985 ;
        RECT 65.325 156.825 65.495 157.015 ;
        RECT 68.085 156.845 68.255 157.035 ;
        RECT 68.545 156.845 68.715 157.035 ;
        RECT 70.385 156.845 70.555 157.035 ;
        RECT 74.525 156.825 74.695 157.015 ;
        RECT 75.440 156.845 75.610 157.035 ;
        RECT 76.365 156.985 76.535 157.015 ;
        RECT 76.365 156.875 76.540 156.985 ;
        RECT 76.365 156.825 76.535 156.875 ;
        RECT 76.830 156.825 77.000 157.015 ;
        RECT 80.040 156.845 80.210 157.035 ;
        RECT 80.510 156.825 80.680 157.015 ;
        RECT 84.645 156.870 84.805 156.980 ;
        RECT 88.325 156.825 88.495 157.015 ;
        RECT 90.165 156.845 90.335 157.035 ;
        RECT 90.680 156.875 90.800 156.985 ;
        RECT 91.545 156.825 91.715 157.015 ;
        RECT 92.465 156.845 92.635 157.035 ;
        RECT 92.925 156.845 93.095 157.035 ;
        RECT 94.360 156.875 94.480 156.985 ;
        RECT 96.145 156.845 96.315 157.035 ;
        RECT 96.605 156.845 96.775 157.035 ;
        RECT 97.065 156.825 97.235 157.015 ;
        RECT 99.365 156.845 99.535 157.035 ;
        RECT 99.825 156.845 99.995 157.035 ;
        RECT 100.740 156.825 100.910 157.015 ;
        RECT 101.260 156.875 101.380 156.985 ;
        RECT 102.180 156.875 102.300 156.985 ;
        RECT 103.045 156.825 103.215 157.015 ;
        RECT 103.510 156.825 103.680 157.015 ;
        RECT 103.965 156.845 104.135 157.035 ;
        RECT 105.345 156.845 105.515 157.035 ;
        RECT 105.805 156.845 105.975 157.035 ;
        RECT 107.645 156.880 107.805 156.990 ;
        RECT 108.110 156.845 108.280 157.035 ;
        RECT 110.400 156.825 110.570 157.015 ;
        RECT 112.245 156.880 112.405 156.990 ;
        RECT 114.085 156.825 114.255 157.015 ;
        RECT 115.925 156.825 116.095 157.035 ;
        RECT 116.385 157.015 116.555 157.035 ;
        RECT 116.385 156.845 116.560 157.015 ;
        RECT 116.390 156.825 116.560 156.845 ;
        RECT 120.525 156.825 120.695 157.015 ;
        RECT 126.045 156.825 126.215 157.035 ;
        RECT 127.425 156.825 127.595 157.035 ;
        RECT 14.585 156.015 15.955 156.825 ;
        RECT 17.255 156.145 26.535 156.825 ;
        RECT 17.255 156.025 19.590 156.145 ;
        RECT 17.255 155.915 18.175 156.025 ;
        RECT 24.255 155.925 25.175 156.145 ;
        RECT 26.545 156.045 27.915 156.825 ;
        RECT 27.925 156.015 29.295 156.825 ;
        RECT 29.305 156.015 32.975 156.825 ;
        RECT 33.215 156.145 37.115 156.825 ;
        RECT 36.185 155.915 37.115 156.145 ;
        RECT 37.135 155.955 37.565 156.740 ;
        RECT 38.045 156.015 39.875 156.825 ;
        RECT 39.885 155.915 43.360 156.825 ;
        RECT 43.565 155.915 47.040 156.825 ;
        RECT 47.245 155.915 50.720 156.825 ;
        RECT 51.385 156.015 53.215 156.825 ;
        RECT 53.595 156.145 62.875 156.825 ;
        RECT 53.595 156.025 55.930 156.145 ;
        RECT 53.595 155.915 54.515 156.025 ;
        RECT 60.595 155.925 61.515 156.145 ;
        RECT 62.895 155.955 63.325 156.740 ;
        RECT 63.805 156.015 65.635 156.825 ;
        RECT 65.730 156.145 74.835 156.825 ;
        RECT 74.845 156.015 76.675 156.825 ;
        RECT 76.685 155.915 80.160 156.825 ;
        RECT 80.365 155.915 83.840 156.825 ;
        RECT 84.965 156.015 88.635 156.825 ;
        RECT 88.655 155.955 89.085 156.740 ;
        RECT 89.105 156.015 91.855 156.825 ;
        RECT 91.865 156.015 97.375 156.825 ;
        RECT 97.580 155.915 101.055 156.825 ;
        RECT 101.525 156.015 103.355 156.825 ;
        RECT 103.365 155.915 106.840 156.825 ;
        RECT 107.240 155.915 110.715 156.825 ;
        RECT 110.725 156.015 114.395 156.825 ;
        RECT 114.415 155.955 114.845 156.740 ;
        RECT 114.865 156.015 116.235 156.825 ;
        RECT 116.245 155.915 118.855 156.825 ;
        RECT 119.005 156.015 120.835 156.825 ;
        RECT 120.845 156.015 126.355 156.825 ;
        RECT 126.365 156.015 127.735 156.825 ;
      LAYER nwell ;
        RECT 14.390 152.795 127.930 155.625 ;
      LAYER pwell ;
        RECT 14.585 151.595 15.955 152.405 ;
        RECT 16.425 151.595 20.095 152.405 ;
        RECT 23.305 152.275 24.235 152.505 ;
        RECT 20.335 151.595 24.235 152.275 ;
        RECT 24.255 151.680 24.685 152.465 ;
        RECT 24.705 151.595 26.075 152.405 ;
        RECT 26.085 151.595 29.755 152.405 ;
        RECT 30.135 152.395 31.055 152.505 ;
        RECT 30.135 152.275 32.470 152.395 ;
        RECT 37.135 152.275 38.055 152.495 ;
        RECT 30.135 151.595 39.415 152.275 ;
        RECT 39.425 151.595 42.900 152.505 ;
        RECT 43.105 151.595 44.475 152.405 ;
        RECT 44.485 151.595 49.995 152.405 ;
        RECT 50.015 151.680 50.445 152.465 ;
        RECT 51.385 151.595 56.895 152.405 ;
        RECT 56.915 151.595 58.265 152.505 ;
        RECT 58.655 152.395 59.575 152.505 ;
        RECT 58.655 152.275 60.990 152.395 ;
        RECT 65.655 152.275 66.575 152.495 ;
        RECT 58.655 151.595 67.935 152.275 ;
        RECT 68.405 151.595 71.155 152.405 ;
        RECT 71.650 152.275 72.995 152.505 ;
        RECT 71.165 151.595 72.995 152.275 ;
        RECT 73.005 151.595 75.725 152.505 ;
        RECT 75.775 151.680 76.205 152.465 ;
        RECT 77.145 151.595 80.815 152.405 ;
        RECT 80.825 151.595 86.335 152.405 ;
        RECT 86.715 152.395 87.635 152.505 ;
        RECT 86.715 152.275 89.050 152.395 ;
        RECT 93.715 152.275 94.635 152.495 ;
        RECT 86.715 151.595 95.995 152.275 ;
        RECT 96.005 151.595 101.515 152.405 ;
        RECT 101.535 151.680 101.965 152.465 ;
        RECT 102.445 152.305 103.390 152.505 ;
        RECT 102.445 151.625 105.195 152.305 ;
        RECT 102.445 151.595 103.390 151.625 ;
        RECT 14.725 151.385 14.895 151.595 ;
        RECT 16.160 151.435 16.280 151.545 ;
        RECT 19.785 151.405 19.955 151.595 ;
        RECT 23.650 151.405 23.820 151.595 ;
        RECT 25.765 151.385 25.935 151.595 ;
        RECT 27.145 151.385 27.315 151.575 ;
        RECT 29.445 151.405 29.615 151.595 ;
        RECT 32.665 151.385 32.835 151.575 ;
        RECT 33.125 151.385 33.295 151.575 ;
        RECT 35.425 151.385 35.595 151.575 ;
        RECT 35.885 151.385 36.055 151.575 ;
        RECT 39.105 151.405 39.275 151.595 ;
        RECT 39.570 151.405 39.740 151.595 ;
        RECT 40.945 151.385 41.115 151.575 ;
        RECT 41.410 151.385 41.580 151.575 ;
        RECT 44.165 151.405 44.335 151.595 ;
        RECT 48.305 151.385 48.475 151.575 ;
        RECT 14.585 150.575 15.955 151.385 ;
        RECT 16.795 150.705 26.075 151.385 ;
        RECT 16.795 150.585 19.130 150.705 ;
        RECT 16.795 150.475 17.715 150.585 ;
        RECT 23.795 150.485 24.715 150.705 ;
        RECT 26.085 150.575 27.455 151.385 ;
        RECT 27.465 150.575 32.975 151.385 ;
        RECT 32.995 150.475 34.345 151.385 ;
        RECT 34.365 150.575 35.735 151.385 ;
        RECT 35.745 150.605 37.115 151.385 ;
        RECT 37.135 150.515 37.565 151.300 ;
        RECT 37.585 150.575 41.255 151.385 ;
        RECT 41.265 150.475 44.740 151.385 ;
        RECT 44.945 150.575 48.615 151.385 ;
        RECT 48.770 151.355 48.940 151.575 ;
        RECT 49.685 151.405 49.855 151.595 ;
        RECT 51.065 151.440 51.225 151.550 ;
        RECT 51.530 151.385 51.700 151.575 ;
        RECT 56.585 151.385 56.755 151.595 ;
        RECT 57.045 151.405 57.215 151.595 ;
        RECT 60.450 151.385 60.620 151.575 ;
        RECT 61.240 151.435 61.360 151.545 ;
        RECT 62.565 151.385 62.735 151.575 ;
        RECT 63.540 151.435 63.660 151.545 ;
        RECT 63.945 151.385 64.115 151.575 ;
        RECT 65.380 151.435 65.500 151.545 ;
        RECT 67.165 151.385 67.335 151.575 ;
        RECT 67.625 151.385 67.795 151.595 ;
        RECT 68.140 151.435 68.260 151.545 ;
        RECT 70.845 151.385 71.015 151.595 ;
        RECT 71.305 151.405 71.475 151.595 ;
        RECT 73.145 151.405 73.315 151.595 ;
        RECT 73.605 151.385 73.775 151.575 ;
        RECT 74.525 151.430 74.685 151.540 ;
        RECT 74.985 151.385 75.155 151.575 ;
        RECT 76.825 151.440 76.985 151.550 ;
        RECT 50.430 151.355 51.375 151.385 ;
        RECT 48.625 150.675 51.375 151.355 ;
        RECT 50.430 150.475 51.375 150.675 ;
        RECT 51.385 150.475 54.860 151.385 ;
        RECT 55.065 150.575 56.895 151.385 ;
        RECT 57.135 150.705 61.035 151.385 ;
        RECT 60.105 150.475 61.035 150.705 ;
        RECT 61.505 150.605 62.875 151.385 ;
        RECT 62.895 150.515 63.325 151.300 ;
        RECT 63.805 150.605 65.175 151.385 ;
        RECT 65.645 150.575 67.475 151.385 ;
        RECT 67.485 150.705 69.315 151.385 ;
        RECT 67.970 150.475 69.315 150.705 ;
        RECT 69.325 150.705 71.155 151.385 ;
        RECT 71.175 150.705 73.915 151.385 ;
        RECT 74.845 150.705 77.585 151.385 ;
        RECT 77.605 151.355 78.550 151.385 ;
        RECT 80.040 151.355 80.210 151.575 ;
        RECT 80.505 151.545 80.675 151.595 ;
        RECT 80.505 151.435 80.680 151.545 ;
        RECT 80.505 151.405 80.675 151.435 ;
        RECT 84.185 151.385 84.355 151.575 ;
        RECT 86.025 151.405 86.195 151.595 ;
        RECT 88.050 151.385 88.220 151.575 ;
        RECT 89.300 151.435 89.420 151.545 ;
        RECT 90.625 151.385 90.795 151.575 ;
        RECT 91.545 151.430 91.705 151.540 ;
        RECT 92.005 151.385 92.175 151.575 ;
        RECT 94.305 151.385 94.475 151.575 ;
        RECT 95.685 151.405 95.855 151.595 ;
        RECT 96.145 151.385 96.315 151.575 ;
        RECT 101.205 151.405 101.375 151.595 ;
        RECT 102.180 151.435 102.300 151.545 ;
        RECT 104.880 151.405 105.050 151.625 ;
        RECT 105.205 151.595 108.680 152.505 ;
        RECT 108.885 151.595 112.360 152.505 ;
        RECT 113.025 151.595 118.535 152.405 ;
        RECT 118.555 151.595 119.905 152.505 ;
        RECT 120.385 151.595 121.755 152.375 ;
        RECT 122.685 151.595 126.355 152.405 ;
        RECT 126.365 151.595 127.735 152.405 ;
        RECT 105.350 151.575 105.520 151.595 ;
        RECT 105.345 151.405 105.520 151.575 ;
        RECT 105.345 151.385 105.515 151.405 ;
        RECT 106.725 151.385 106.895 151.575 ;
        RECT 107.190 151.385 107.360 151.575 ;
        RECT 109.030 151.405 109.200 151.595 ;
        RECT 110.865 151.385 111.035 151.575 ;
        RECT 112.760 151.435 112.880 151.545 ;
        RECT 115.465 151.430 115.625 151.540 ;
        RECT 118.225 151.405 118.395 151.595 ;
        RECT 119.605 151.405 119.775 151.595 ;
        RECT 120.120 151.435 120.240 151.545 ;
        RECT 120.525 151.405 120.695 151.595 ;
        RECT 122.365 151.440 122.525 151.550 ;
        RECT 124.665 151.385 124.835 151.575 ;
        RECT 126.045 151.385 126.215 151.595 ;
        RECT 127.425 151.385 127.595 151.595 ;
        RECT 69.325 150.475 70.670 150.705 ;
        RECT 77.605 150.675 80.355 151.355 ;
        RECT 77.605 150.475 78.550 150.675 ;
        RECT 80.825 150.575 84.495 151.385 ;
        RECT 84.735 150.705 88.635 151.385 ;
        RECT 87.705 150.475 88.635 150.705 ;
        RECT 88.655 150.515 89.085 151.300 ;
        RECT 89.575 150.475 90.925 151.385 ;
        RECT 91.865 150.605 93.235 151.385 ;
        RECT 93.255 150.475 94.605 151.385 ;
        RECT 94.625 150.575 96.455 151.385 ;
        RECT 96.465 150.705 105.655 151.385 ;
        RECT 96.465 150.475 97.385 150.705 ;
        RECT 100.215 150.485 101.145 150.705 ;
        RECT 105.665 150.575 107.035 151.385 ;
        RECT 107.045 150.475 110.520 151.385 ;
        RECT 110.835 150.705 114.300 151.385 ;
        RECT 113.380 150.475 114.300 150.705 ;
        RECT 114.415 150.515 114.845 151.300 ;
        RECT 115.785 150.705 124.975 151.385 ;
        RECT 115.785 150.475 116.705 150.705 ;
        RECT 119.535 150.485 120.465 150.705 ;
        RECT 124.985 150.575 126.355 151.385 ;
        RECT 126.365 150.575 127.735 151.385 ;
      LAYER nwell ;
        RECT 14.390 147.355 127.930 150.185 ;
      LAYER pwell ;
        RECT 14.585 146.155 15.955 146.965 ;
        RECT 16.425 146.155 20.095 146.965 ;
        RECT 23.305 146.835 24.235 147.065 ;
        RECT 20.335 146.155 24.235 146.835 ;
        RECT 24.255 146.240 24.685 147.025 ;
        RECT 24.705 146.155 26.075 146.935 ;
        RECT 26.085 146.155 27.915 146.965 ;
        RECT 27.925 146.155 29.295 146.935 ;
        RECT 29.305 146.835 30.235 147.065 ;
        RECT 29.305 146.155 33.205 146.835 ;
        RECT 33.905 146.155 35.735 146.965 ;
        RECT 35.940 146.155 39.415 147.065 ;
        RECT 39.425 146.155 42.900 147.065 ;
        RECT 43.565 146.155 47.235 146.965 ;
        RECT 49.050 146.865 49.995 147.065 ;
        RECT 47.245 146.185 49.995 146.865 ;
        RECT 50.015 146.240 50.445 147.025 ;
        RECT 14.725 145.945 14.895 146.155 ;
        RECT 16.160 145.995 16.280 146.105 ;
        RECT 19.325 145.945 19.495 146.135 ;
        RECT 19.785 145.945 19.955 146.155 ;
        RECT 21.165 145.945 21.335 146.135 ;
        RECT 23.650 145.965 23.820 146.155 ;
        RECT 25.765 145.965 25.935 146.155 ;
        RECT 27.605 145.965 27.775 146.155 ;
        RECT 28.065 145.965 28.235 146.155 ;
        RECT 29.720 145.965 29.890 146.155 ;
        RECT 31.745 145.945 31.915 146.135 ;
        RECT 33.125 145.945 33.295 146.135 ;
        RECT 33.640 145.995 33.760 146.105 ;
        RECT 35.425 145.965 35.595 146.155 ;
        RECT 36.805 145.945 36.975 146.135 ;
        RECT 37.780 145.995 37.900 146.105 ;
        RECT 39.100 145.965 39.270 146.155 ;
        RECT 39.570 145.965 39.740 146.155 ;
        RECT 40.485 145.945 40.655 146.135 ;
        RECT 40.945 145.945 41.115 146.135 ;
        RECT 43.300 145.995 43.420 146.105 ;
        RECT 46.925 145.965 47.095 146.155 ;
        RECT 47.390 145.965 47.560 146.185 ;
        RECT 49.050 146.155 49.995 146.185 ;
        RECT 50.925 146.155 52.295 146.935 ;
        RECT 53.225 146.155 56.700 147.065 ;
        RECT 56.905 146.155 59.655 146.965 ;
        RECT 62.865 146.835 63.795 147.065 ;
        RECT 59.895 146.155 63.795 146.835 ;
        RECT 63.805 146.155 65.175 146.965 ;
        RECT 65.185 146.155 70.695 146.965 ;
        RECT 70.705 146.835 72.050 147.065 ;
        RECT 73.030 146.835 74.375 147.065 ;
        RECT 70.705 146.155 72.535 146.835 ;
        RECT 72.545 146.155 74.375 146.835 ;
        RECT 74.385 146.155 75.755 146.965 ;
        RECT 75.775 146.240 76.205 147.025 ;
        RECT 76.420 146.155 79.895 147.065 ;
        RECT 79.905 146.155 83.380 147.065 ;
        RECT 83.585 146.155 84.955 146.965 ;
        RECT 85.335 146.955 86.255 147.065 ;
        RECT 85.335 146.835 87.670 146.955 ;
        RECT 92.335 146.835 93.255 147.055 ;
        RECT 85.335 146.155 94.615 146.835 ;
        RECT 95.095 146.155 96.445 147.065 ;
        RECT 99.665 146.835 100.595 147.065 ;
        RECT 96.695 146.155 100.595 146.835 ;
        RECT 101.535 146.240 101.965 147.025 ;
        RECT 101.985 146.155 103.355 146.935 ;
        RECT 103.825 146.865 104.770 147.065 ;
        RECT 103.825 146.185 106.575 146.865 ;
        RECT 103.825 146.155 104.770 146.185 ;
        RECT 50.660 145.995 50.780 146.105 ;
        RECT 51.525 145.945 51.695 146.135 ;
        RECT 51.985 145.965 52.155 146.155 ;
        RECT 52.260 145.945 52.430 146.135 ;
        RECT 52.905 146.000 53.065 146.110 ;
        RECT 53.370 145.965 53.540 146.155 ;
        RECT 56.180 145.995 56.300 146.105 ;
        RECT 57.965 145.945 58.135 146.135 ;
        RECT 58.425 145.945 58.595 146.135 ;
        RECT 59.345 145.965 59.515 146.155 ;
        RECT 59.860 145.995 59.980 146.105 ;
        RECT 62.565 145.945 62.735 146.135 ;
        RECT 63.210 145.965 63.380 146.155 ;
        RECT 63.540 145.995 63.660 146.105 ;
        RECT 64.865 145.965 65.035 146.155 ;
        RECT 67.350 145.945 67.520 146.135 ;
        RECT 68.140 145.995 68.260 146.105 ;
        RECT 70.385 145.965 70.555 146.155 ;
        RECT 72.225 145.965 72.395 146.155 ;
        RECT 72.685 145.965 72.855 146.155 ;
        RECT 73.605 145.945 73.775 146.135 ;
        RECT 75.445 145.965 75.615 146.155 ;
        RECT 79.580 146.135 79.750 146.155 ;
        RECT 79.125 145.945 79.295 146.135 ;
        RECT 79.580 145.965 79.760 146.135 ;
        RECT 80.050 145.965 80.220 146.155 ;
        RECT 82.400 145.995 82.520 146.105 ;
        RECT 14.585 145.135 15.955 145.945 ;
        RECT 15.965 145.135 19.635 145.945 ;
        RECT 19.655 145.035 21.005 145.945 ;
        RECT 21.035 145.035 22.385 145.945 ;
        RECT 22.775 145.265 32.055 145.945 ;
        RECT 22.775 145.145 25.110 145.265 ;
        RECT 22.775 145.035 23.695 145.145 ;
        RECT 29.775 145.045 30.695 145.265 ;
        RECT 32.065 145.135 33.435 145.945 ;
        RECT 33.445 145.135 37.115 145.945 ;
        RECT 37.135 145.075 37.565 145.860 ;
        RECT 38.045 145.135 40.795 145.945 ;
        RECT 40.815 145.035 42.165 145.945 ;
        RECT 42.555 145.265 51.835 145.945 ;
        RECT 51.845 145.265 55.745 145.945 ;
        RECT 42.555 145.145 44.890 145.265 ;
        RECT 42.555 145.035 43.475 145.145 ;
        RECT 49.555 145.045 50.475 145.265 ;
        RECT 51.845 145.035 52.775 145.265 ;
        RECT 56.445 145.135 58.275 145.945 ;
        RECT 58.295 145.035 59.645 145.945 ;
        RECT 60.125 145.135 62.875 145.945 ;
        RECT 62.895 145.075 63.325 145.860 ;
        RECT 64.035 145.265 67.935 145.945 ;
        RECT 67.005 145.035 67.935 145.265 ;
        RECT 68.405 145.135 73.915 145.945 ;
        RECT 73.925 145.135 79.435 145.945 ;
        RECT 79.590 145.915 79.760 145.965 ;
        RECT 84.185 145.945 84.355 146.135 ;
        RECT 84.645 145.965 84.815 146.155 ;
        RECT 88.050 145.945 88.220 146.135 ;
        RECT 89.705 145.990 89.865 146.100 ;
        RECT 90.165 145.945 90.335 146.135 ;
        RECT 91.600 145.995 91.720 146.105 ;
        RECT 93.385 145.945 93.555 146.135 ;
        RECT 93.845 145.945 94.015 146.135 ;
        RECT 94.305 145.965 94.475 146.155 ;
        RECT 94.820 145.995 94.940 146.105 ;
        RECT 95.225 145.965 95.395 146.155 ;
        RECT 97.580 145.995 97.700 146.105 ;
        RECT 100.010 145.965 100.180 146.155 ;
        RECT 101.205 145.945 101.375 146.135 ;
        RECT 102.125 145.965 102.295 146.155 ;
        RECT 103.560 145.995 103.680 146.105 ;
        RECT 106.260 145.965 106.430 146.185 ;
        RECT 106.585 146.155 110.060 147.065 ;
        RECT 110.265 146.155 112.095 146.965 ;
        RECT 115.305 146.835 116.235 147.065 ;
        RECT 112.335 146.155 116.235 146.835 ;
        RECT 116.615 146.955 117.535 147.065 ;
        RECT 116.615 146.835 118.950 146.955 ;
        RECT 123.615 146.835 124.535 147.055 ;
        RECT 116.615 146.155 125.895 146.835 ;
        RECT 126.365 146.155 127.735 146.965 ;
        RECT 106.730 146.135 106.900 146.155 ;
        RECT 106.725 145.965 106.900 146.135 ;
        RECT 106.725 145.945 106.895 145.965 ;
        RECT 81.250 145.915 82.195 145.945 ;
        RECT 79.445 145.235 82.195 145.915 ;
        RECT 81.250 145.035 82.195 145.235 ;
        RECT 82.665 145.135 84.495 145.945 ;
        RECT 84.735 145.265 88.635 145.945 ;
        RECT 87.705 145.035 88.635 145.265 ;
        RECT 88.655 145.075 89.085 145.860 ;
        RECT 90.025 145.165 91.395 145.945 ;
        RECT 91.865 145.135 93.695 145.945 ;
        RECT 93.815 145.265 97.280 145.945 ;
        RECT 96.360 145.035 97.280 145.265 ;
        RECT 97.845 145.135 101.515 145.945 ;
        RECT 101.525 145.135 107.035 145.945 ;
        RECT 107.190 145.915 107.360 146.135 ;
        RECT 109.950 145.945 110.120 146.135 ;
        RECT 111.785 145.965 111.955 146.155 ;
        RECT 114.085 145.990 114.245 146.100 ;
        RECT 115.060 145.995 115.180 146.105 ;
        RECT 115.650 145.965 115.820 146.155 ;
        RECT 118.870 145.945 119.040 146.135 ;
        RECT 119.605 145.945 119.775 146.135 ;
        RECT 121.040 145.995 121.160 146.105 ;
        RECT 121.445 145.945 121.615 146.135 ;
        RECT 125.585 145.965 125.755 146.155 ;
        RECT 126.045 146.105 126.215 146.135 ;
        RECT 126.045 145.995 126.220 146.105 ;
        RECT 126.045 145.945 126.215 145.995 ;
        RECT 127.425 145.945 127.595 146.155 ;
        RECT 108.850 145.915 109.795 145.945 ;
        RECT 107.045 145.235 109.795 145.915 ;
        RECT 108.850 145.035 109.795 145.235 ;
        RECT 109.805 145.035 113.280 145.945 ;
        RECT 114.415 145.075 114.845 145.860 ;
        RECT 115.555 145.265 119.455 145.945 ;
        RECT 118.525 145.035 119.455 145.265 ;
        RECT 119.475 145.035 120.825 145.945 ;
        RECT 121.305 145.165 122.675 145.945 ;
        RECT 122.685 145.135 126.355 145.945 ;
        RECT 126.365 145.135 127.735 145.945 ;
      LAYER nwell ;
        RECT 14.390 141.915 127.930 144.745 ;
      LAYER pwell ;
        RECT 14.585 140.715 15.955 141.525 ;
        RECT 15.965 140.715 18.715 141.525 ;
        RECT 18.725 140.715 24.235 141.525 ;
        RECT 24.255 140.800 24.685 141.585 ;
        RECT 25.165 140.715 28.835 141.525 ;
        RECT 28.845 140.715 34.355 141.525 ;
        RECT 34.365 141.425 35.310 141.625 ;
        RECT 34.365 140.745 37.115 141.425 ;
        RECT 34.365 140.715 35.310 140.745 ;
        RECT 14.725 140.505 14.895 140.715 ;
        RECT 18.405 140.525 18.575 140.715 ;
        RECT 23.925 140.525 24.095 140.715 ;
        RECT 24.900 140.555 25.020 140.665 ;
        RECT 25.305 140.505 25.475 140.695 ;
        RECT 28.065 140.505 28.235 140.695 ;
        RECT 28.525 140.525 28.695 140.715 ;
        RECT 33.585 140.505 33.755 140.695 ;
        RECT 34.045 140.525 34.215 140.715 ;
        RECT 36.800 140.525 36.970 140.745 ;
        RECT 38.045 140.715 41.715 141.525 ;
        RECT 41.725 140.715 47.235 141.525 ;
        RECT 47.245 141.425 48.190 141.625 ;
        RECT 47.245 140.745 49.995 141.425 ;
        RECT 50.015 140.800 50.445 141.585 ;
        RECT 47.245 140.715 48.190 140.745 ;
        RECT 37.725 140.560 37.885 140.670 ;
        RECT 38.185 140.550 38.345 140.660 ;
        RECT 34.065 140.505 34.215 140.525 ;
        RECT 14.585 139.695 15.955 140.505 ;
        RECT 16.335 139.825 25.615 140.505 ;
        RECT 16.335 139.705 18.670 139.825 ;
        RECT 16.335 139.595 17.255 139.705 ;
        RECT 23.335 139.605 24.255 139.825 ;
        RECT 25.625 139.695 28.375 140.505 ;
        RECT 28.385 139.695 33.895 140.505 ;
        RECT 34.065 139.685 35.995 140.505 ;
        RECT 38.505 140.475 39.450 140.505 ;
        RECT 40.940 140.475 41.110 140.695 ;
        RECT 41.405 140.665 41.575 140.715 ;
        RECT 41.405 140.555 41.580 140.665 ;
        RECT 41.405 140.525 41.575 140.555 ;
        RECT 44.165 140.505 44.335 140.695 ;
        RECT 46.925 140.525 47.095 140.715 ;
        RECT 49.680 140.695 49.850 140.745 ;
        RECT 50.465 140.715 52.295 141.525 ;
        RECT 52.305 140.715 55.780 141.625 ;
        RECT 58.640 141.395 59.560 141.625 ;
        RECT 56.095 140.715 59.560 141.395 ;
        RECT 59.665 141.395 60.585 141.625 ;
        RECT 63.415 141.395 64.345 141.615 ;
        RECT 59.665 140.715 68.855 141.395 ;
        RECT 68.865 140.715 70.235 141.495 ;
        RECT 70.245 140.715 71.615 141.525 ;
        RECT 71.635 140.715 72.985 141.625 ;
        RECT 73.005 140.715 75.755 141.525 ;
        RECT 75.775 140.800 76.205 141.585 ;
        RECT 76.685 140.715 79.435 141.525 ;
        RECT 79.445 140.715 84.955 141.525 ;
        RECT 84.965 140.715 90.475 141.525 ;
        RECT 90.485 140.715 95.995 141.525 ;
        RECT 96.005 140.715 101.515 141.525 ;
        RECT 101.535 140.800 101.965 141.585 ;
        RECT 101.985 140.715 104.735 141.525 ;
        RECT 104.745 140.715 110.255 141.525 ;
        RECT 110.265 140.715 115.775 141.525 ;
        RECT 118.985 141.395 119.915 141.625 ;
        RECT 116.015 140.715 119.915 141.395 ;
        RECT 119.935 140.715 121.285 141.625 ;
        RECT 121.305 140.715 122.675 141.525 ;
        RECT 122.685 140.715 126.355 141.525 ;
        RECT 126.365 140.715 127.735 141.525 ;
        RECT 49.680 140.525 49.855 140.695 ;
        RECT 51.985 140.525 52.155 140.715 ;
        RECT 52.450 140.525 52.620 140.715 ;
        RECT 49.685 140.505 49.855 140.525 ;
        RECT 55.205 140.505 55.375 140.695 ;
        RECT 55.665 140.505 55.835 140.695 ;
        RECT 56.125 140.525 56.295 140.715 ;
        RECT 57.100 140.555 57.220 140.665 ;
        RECT 58.885 140.505 59.055 140.695 ;
        RECT 59.350 140.505 59.520 140.695 ;
        RECT 63.540 140.555 63.660 140.665 ;
        RECT 63.950 140.505 64.120 140.695 ;
        RECT 68.545 140.525 68.715 140.715 ;
        RECT 69.925 140.525 70.095 140.715 ;
        RECT 71.305 140.525 71.475 140.715 ;
        RECT 72.685 140.525 72.855 140.715 ;
        RECT 75.445 140.525 75.615 140.715 ;
        RECT 76.420 140.555 76.540 140.665 ;
        RECT 76.825 140.505 76.995 140.695 ;
        RECT 77.340 140.555 77.460 140.665 ;
        RECT 79.125 140.505 79.295 140.715 ;
        RECT 79.590 140.505 79.760 140.695 ;
        RECT 84.185 140.505 84.355 140.695 ;
        RECT 84.645 140.525 84.815 140.715 ;
        RECT 88.050 140.505 88.220 140.695 ;
        RECT 89.245 140.505 89.415 140.695 ;
        RECT 90.165 140.525 90.335 140.715 ;
        RECT 92.005 140.505 92.175 140.695 ;
        RECT 95.685 140.525 95.855 140.715 ;
        RECT 97.525 140.505 97.695 140.695 ;
        RECT 101.205 140.525 101.375 140.715 ;
        RECT 104.425 140.525 104.595 140.715 ;
        RECT 107.185 140.505 107.355 140.695 ;
        RECT 107.700 140.555 107.820 140.665 ;
        RECT 109.485 140.505 109.655 140.695 ;
        RECT 109.945 140.525 110.115 140.715 ;
        RECT 113.160 140.505 113.330 140.695 ;
        RECT 114.085 140.550 114.245 140.660 ;
        RECT 115.060 140.555 115.180 140.665 ;
        RECT 115.465 140.505 115.635 140.715 ;
        RECT 119.330 140.525 119.500 140.715 ;
        RECT 120.065 140.525 120.235 140.715 ;
        RECT 122.365 140.525 122.535 140.715 ;
        RECT 126.045 140.505 126.215 140.715 ;
        RECT 127.425 140.505 127.595 140.715 ;
        RECT 35.045 139.595 35.995 139.685 ;
        RECT 37.135 139.635 37.565 140.420 ;
        RECT 38.505 139.795 41.255 140.475 ;
        RECT 38.505 139.595 39.450 139.795 ;
        RECT 41.725 139.695 44.475 140.505 ;
        RECT 44.485 139.695 49.995 140.505 ;
        RECT 50.005 139.695 55.515 140.505 ;
        RECT 55.535 139.595 56.885 140.505 ;
        RECT 57.365 139.695 59.195 140.505 ;
        RECT 59.205 139.595 62.680 140.505 ;
        RECT 62.895 139.635 63.325 140.420 ;
        RECT 63.805 139.595 67.280 140.505 ;
        RECT 67.855 139.825 77.135 140.505 ;
        RECT 67.855 139.705 70.190 139.825 ;
        RECT 67.855 139.595 68.775 139.705 ;
        RECT 74.855 139.605 75.775 139.825 ;
        RECT 77.605 139.695 79.435 140.505 ;
        RECT 79.445 139.595 82.920 140.505 ;
        RECT 83.125 139.695 84.495 140.505 ;
        RECT 84.735 139.825 88.635 140.505 ;
        RECT 87.705 139.595 88.635 139.825 ;
        RECT 88.655 139.635 89.085 140.420 ;
        RECT 89.105 139.725 90.475 140.505 ;
        RECT 90.485 139.695 92.315 140.505 ;
        RECT 92.325 139.695 97.835 140.505 ;
        RECT 98.215 139.825 107.495 140.505 ;
        RECT 98.215 139.705 100.550 139.825 ;
        RECT 98.215 139.595 99.135 139.705 ;
        RECT 105.215 139.605 106.135 139.825 ;
        RECT 107.965 139.695 109.795 140.505 ;
        RECT 110.000 139.595 113.475 140.505 ;
        RECT 114.415 139.635 114.845 140.420 ;
        RECT 115.335 139.595 116.685 140.505 ;
        RECT 117.075 139.825 126.355 140.505 ;
        RECT 117.075 139.705 119.410 139.825 ;
        RECT 117.075 139.595 117.995 139.705 ;
        RECT 124.075 139.605 124.995 139.825 ;
        RECT 126.365 139.695 127.735 140.505 ;
      LAYER nwell ;
        RECT 14.390 136.475 127.930 139.305 ;
      LAYER pwell ;
        RECT 14.585 135.275 15.955 136.085 ;
        RECT 16.425 135.275 20.095 136.085 ;
        RECT 20.105 135.955 21.035 136.185 ;
        RECT 20.105 135.275 24.005 135.955 ;
        RECT 24.255 135.360 24.685 136.145 ;
        RECT 24.705 135.275 28.375 136.085 ;
        RECT 28.385 135.955 29.315 136.185 ;
        RECT 33.665 136.095 34.615 136.185 ;
        RECT 28.385 135.275 32.285 135.955 ;
        RECT 32.685 135.275 34.615 136.095 ;
        RECT 34.825 135.985 35.770 136.185 ;
        RECT 37.585 135.985 38.530 136.185 ;
        RECT 34.825 135.305 37.575 135.985 ;
        RECT 37.585 135.305 40.335 135.985 ;
        RECT 34.825 135.275 35.770 135.305 ;
        RECT 14.725 135.065 14.895 135.275 ;
        RECT 16.160 135.115 16.280 135.225 ;
        RECT 17.485 135.065 17.655 135.255 ;
        RECT 17.945 135.065 18.115 135.255 ;
        RECT 19.325 135.065 19.495 135.255 ;
        RECT 19.785 135.085 19.955 135.275 ;
        RECT 20.520 135.085 20.690 135.275 ;
        RECT 28.065 135.085 28.235 135.275 ;
        RECT 28.800 135.085 28.970 135.275 ;
        RECT 32.685 135.255 32.835 135.275 ;
        RECT 29.905 135.065 30.075 135.255 ;
        RECT 30.420 135.115 30.540 135.225 ;
        RECT 30.825 135.085 30.995 135.255 ;
        RECT 32.665 135.085 32.835 135.255 ;
        RECT 30.845 135.065 30.995 135.085 ;
        RECT 36.530 135.065 36.700 135.255 ;
        RECT 37.260 135.085 37.430 135.305 ;
        RECT 37.585 135.275 38.530 135.305 ;
        RECT 39.105 135.065 39.275 135.255 ;
        RECT 14.585 134.255 15.955 135.065 ;
        RECT 16.435 134.155 17.785 135.065 ;
        RECT 17.805 134.285 19.175 135.065 ;
        RECT 19.195 134.155 20.545 135.065 ;
        RECT 20.935 134.385 30.215 135.065 ;
        RECT 20.935 134.265 23.270 134.385 ;
        RECT 20.935 134.155 21.855 134.265 ;
        RECT 27.935 134.165 28.855 134.385 ;
        RECT 30.845 134.245 32.775 135.065 ;
        RECT 33.215 134.385 37.115 135.065 ;
        RECT 31.825 134.155 32.775 134.245 ;
        RECT 36.185 134.155 37.115 134.385 ;
        RECT 37.135 134.195 37.565 134.980 ;
        RECT 37.585 134.255 39.415 135.065 ;
        RECT 39.570 135.035 39.740 135.255 ;
        RECT 40.020 135.085 40.190 135.305 ;
        RECT 40.805 135.275 43.555 136.085 ;
        RECT 43.565 135.985 44.510 136.185 ;
        RECT 43.565 135.305 46.315 135.985 ;
        RECT 43.565 135.275 44.510 135.305 ;
        RECT 40.540 135.115 40.660 135.225 ;
        RECT 41.230 135.035 42.175 135.065 ;
        RECT 42.330 135.035 42.500 135.255 ;
        RECT 43.245 135.085 43.415 135.275 ;
        RECT 45.090 135.065 45.260 135.255 ;
        RECT 46.000 135.085 46.170 135.305 ;
        RECT 46.325 135.275 49.800 136.185 ;
        RECT 50.015 135.360 50.445 136.145 ;
        RECT 50.465 135.275 53.215 136.085 ;
        RECT 56.425 135.955 57.355 136.185 ;
        RECT 53.455 135.275 57.355 135.955 ;
        RECT 57.825 135.275 59.195 136.055 ;
        RECT 59.205 135.275 61.035 136.085 ;
        RECT 61.045 135.275 64.520 136.185 ;
        RECT 67.380 135.955 68.300 136.185 ;
        RECT 64.835 135.275 68.300 135.955 ;
        RECT 68.405 135.275 71.615 136.185 ;
        RECT 72.085 135.275 75.755 136.085 ;
        RECT 75.775 135.360 76.205 136.145 ;
        RECT 77.145 135.985 78.090 136.185 ;
        RECT 77.145 135.305 79.895 135.985 ;
        RECT 77.145 135.275 78.090 135.305 ;
        RECT 46.470 135.085 46.640 135.275 ;
        RECT 48.770 135.065 48.940 135.255 ;
        RECT 52.905 135.085 53.075 135.275 ;
        RECT 56.770 135.085 56.940 135.275 ;
        RECT 57.560 135.115 57.680 135.225 ;
        RECT 57.965 135.085 58.135 135.275 ;
        RECT 60.725 135.085 60.895 135.275 ;
        RECT 61.190 135.085 61.360 135.275 ;
        RECT 61.645 135.065 61.815 135.255 ;
        RECT 62.565 135.110 62.725 135.220 ;
        RECT 63.490 135.065 63.660 135.255 ;
        RECT 64.865 135.085 65.035 135.275 ;
        RECT 67.625 135.110 67.785 135.220 ;
        RECT 68.545 135.085 68.715 135.275 ;
        RECT 71.820 135.115 71.940 135.225 ;
        RECT 73.145 135.065 73.315 135.255 ;
        RECT 75.445 135.085 75.615 135.275 ;
        RECT 76.825 135.120 76.985 135.230 ;
        RECT 78.665 135.065 78.835 135.255 ;
        RECT 43.990 135.035 44.935 135.065 ;
        RECT 39.425 134.355 42.175 135.035 ;
        RECT 42.185 134.355 44.935 135.035 ;
        RECT 41.230 134.155 42.175 134.355 ;
        RECT 43.990 134.155 44.935 134.355 ;
        RECT 44.945 134.155 48.420 135.065 ;
        RECT 48.625 134.155 52.100 135.065 ;
        RECT 52.675 134.385 61.955 135.065 ;
        RECT 52.675 134.265 55.010 134.385 ;
        RECT 52.675 134.155 53.595 134.265 ;
        RECT 59.675 134.165 60.595 134.385 ;
        RECT 62.895 134.195 63.325 134.980 ;
        RECT 63.345 134.155 66.820 135.065 ;
        RECT 67.945 134.255 73.455 135.065 ;
        RECT 73.465 134.255 78.975 135.065 ;
        RECT 79.130 135.035 79.300 135.255 ;
        RECT 79.580 135.085 79.750 135.305 ;
        RECT 79.905 135.275 83.380 136.185 ;
        RECT 83.955 136.075 84.875 136.185 ;
        RECT 83.955 135.955 86.290 136.075 ;
        RECT 90.955 135.955 91.875 136.175 ;
        RECT 93.245 135.955 94.175 136.185 ;
        RECT 83.955 135.275 93.235 135.955 ;
        RECT 93.245 135.275 97.145 135.955 ;
        RECT 98.040 135.275 101.515 136.185 ;
        RECT 101.535 135.360 101.965 136.145 ;
        RECT 106.105 135.955 107.035 136.185 ;
        RECT 103.135 135.275 107.035 135.955 ;
        RECT 107.045 135.275 108.415 136.055 ;
        RECT 112.545 135.955 113.475 136.185 ;
        RECT 109.575 135.275 113.475 135.955 ;
        RECT 113.855 136.075 114.775 136.185 ;
        RECT 113.855 135.955 116.190 136.075 ;
        RECT 120.855 135.955 121.775 136.175 ;
        RECT 113.855 135.275 123.135 135.955 ;
        RECT 123.145 135.275 124.515 136.055 ;
        RECT 124.525 135.275 126.355 136.085 ;
        RECT 126.365 135.275 127.735 136.085 ;
        RECT 80.050 135.085 80.220 135.275 ;
        RECT 86.945 135.065 87.115 135.255 ;
        RECT 88.325 135.065 88.495 135.255 ;
        RECT 92.925 135.085 93.095 135.275 ;
        RECT 93.660 135.085 93.830 135.275 ;
        RECT 97.580 135.115 97.700 135.225 ;
        RECT 98.445 135.065 98.615 135.255 ;
        RECT 80.790 135.035 81.735 135.065 ;
        RECT 78.985 134.355 81.735 135.035 ;
        RECT 80.790 134.155 81.735 134.355 ;
        RECT 81.745 134.255 87.255 135.065 ;
        RECT 87.275 134.155 88.625 135.065 ;
        RECT 88.655 134.195 89.085 134.980 ;
        RECT 89.475 134.385 98.755 135.065 ;
        RECT 98.765 135.035 99.710 135.065 ;
        RECT 101.200 135.035 101.370 135.275 ;
        RECT 102.585 135.065 102.755 135.255 ;
        RECT 103.100 135.115 103.220 135.225 ;
        RECT 89.475 134.265 91.810 134.385 ;
        RECT 89.475 134.155 90.395 134.265 ;
        RECT 96.475 134.165 97.395 134.385 ;
        RECT 98.765 134.355 101.515 135.035 ;
        RECT 98.765 134.155 99.710 134.355 ;
        RECT 101.535 134.155 102.885 135.065 ;
        RECT 103.365 135.035 104.310 135.065 ;
        RECT 105.800 135.035 105.970 135.255 ;
        RECT 106.270 135.065 106.440 135.255 ;
        RECT 106.450 135.085 106.620 135.275 ;
        RECT 108.105 135.085 108.275 135.275 ;
        RECT 109.025 135.120 109.185 135.230 ;
        RECT 103.365 134.355 106.115 135.035 ;
        RECT 103.365 134.155 104.310 134.355 ;
        RECT 106.125 134.155 109.600 135.065 ;
        RECT 109.805 135.035 110.750 135.065 ;
        RECT 112.240 135.035 112.410 135.255 ;
        RECT 112.890 135.085 113.060 135.275 ;
        RECT 114.085 135.065 114.255 135.255 ;
        RECT 115.060 135.115 115.180 135.225 ;
        RECT 118.685 135.065 118.855 135.255 ;
        RECT 119.145 135.065 119.315 135.255 ;
        RECT 120.580 135.115 120.700 135.225 ;
        RECT 122.825 135.085 122.995 135.275 ;
        RECT 123.285 135.085 123.455 135.275 ;
        RECT 126.045 135.065 126.215 135.275 ;
        RECT 127.425 135.065 127.595 135.275 ;
        RECT 109.805 134.355 112.555 135.035 ;
        RECT 109.805 134.155 110.750 134.355 ;
        RECT 112.565 134.255 114.395 135.065 ;
        RECT 114.415 134.195 114.845 134.980 ;
        RECT 115.325 134.255 118.995 135.065 ;
        RECT 119.005 134.285 120.375 135.065 ;
        RECT 120.845 134.255 126.355 135.065 ;
        RECT 126.365 134.255 127.735 135.065 ;
      LAYER nwell ;
        RECT 14.390 131.035 127.930 133.865 ;
      LAYER pwell ;
        RECT 14.585 129.835 15.955 130.645 ;
        RECT 16.425 129.835 20.095 130.645 ;
        RECT 23.305 130.515 24.235 130.745 ;
        RECT 20.335 129.835 24.235 130.515 ;
        RECT 24.255 129.920 24.685 130.705 ;
        RECT 25.165 129.835 28.835 130.645 ;
        RECT 30.595 130.635 31.515 130.745 ;
        RECT 28.845 129.835 30.215 130.615 ;
        RECT 30.595 130.515 32.930 130.635 ;
        RECT 37.595 130.515 38.515 130.735 ;
        RECT 30.595 129.835 39.875 130.515 ;
        RECT 39.970 129.835 49.075 130.515 ;
        RECT 50.015 129.920 50.445 130.705 ;
        RECT 50.925 129.835 54.595 130.645 ;
        RECT 54.605 129.835 60.115 130.645 ;
        RECT 60.125 129.835 65.635 130.645 ;
        RECT 68.845 130.515 69.775 130.745 ;
        RECT 71.825 130.655 72.775 130.745 ;
        RECT 65.875 129.835 69.775 130.515 ;
        RECT 69.785 129.835 71.615 130.515 ;
        RECT 71.825 129.835 73.755 130.655 ;
        RECT 73.925 129.835 75.755 130.515 ;
        RECT 75.775 129.920 76.205 130.705 ;
        RECT 78.725 130.655 79.675 130.745 ;
        RECT 76.685 129.835 78.515 130.645 ;
        RECT 78.725 129.835 80.655 130.655 ;
        RECT 80.825 129.835 83.575 130.645 ;
        RECT 83.585 129.835 89.095 130.645 ;
        RECT 89.115 129.835 90.465 130.745 ;
        RECT 90.505 129.835 101.515 130.745 ;
        RECT 101.535 129.920 101.965 130.705 ;
        RECT 110.005 130.655 110.955 130.745 ;
        RECT 102.445 129.835 104.275 130.645 ;
        RECT 104.285 129.835 109.795 130.645 ;
        RECT 110.005 129.835 111.935 130.655 ;
        RECT 112.565 129.835 115.315 130.645 ;
        RECT 115.325 129.835 120.835 130.645 ;
        RECT 120.845 129.835 126.355 130.645 ;
        RECT 126.365 129.835 127.735 130.645 ;
        RECT 14.725 129.625 14.895 129.835 ;
        RECT 16.160 129.675 16.280 129.785 ;
        RECT 17.025 129.625 17.195 129.815 ;
        RECT 19.785 129.645 19.955 129.835 ;
        RECT 23.650 129.645 23.820 129.835 ;
        RECT 24.900 129.675 25.020 129.785 ;
        RECT 26.685 129.625 26.855 129.815 ;
        RECT 27.605 129.670 27.765 129.780 ;
        RECT 28.525 129.645 28.695 129.835 ;
        RECT 29.905 129.645 30.075 129.835 ;
        RECT 33.125 129.625 33.295 129.815 ;
        RECT 33.585 129.625 33.755 129.815 ;
        RECT 35.020 129.675 35.140 129.785 ;
        RECT 36.805 129.625 36.975 129.815 ;
        RECT 38.185 129.670 38.345 129.780 ;
        RECT 39.565 129.625 39.735 129.835 ;
        RECT 40.025 129.645 40.195 129.815 ;
        RECT 42.325 129.645 42.495 129.815 ;
        RECT 40.045 129.625 40.195 129.645 ;
        RECT 42.345 129.625 42.495 129.645 ;
        RECT 46.925 129.625 47.095 129.815 ;
        RECT 47.385 129.645 47.555 129.815 ;
        RECT 48.765 129.645 48.935 129.835 ;
        RECT 49.685 129.680 49.845 129.790 ;
        RECT 50.605 129.785 50.775 129.815 ;
        RECT 50.605 129.675 50.780 129.785 ;
        RECT 47.405 129.625 47.555 129.645 ;
        RECT 50.605 129.625 50.775 129.675 ;
        RECT 54.285 129.625 54.455 129.835 ;
        RECT 58.150 129.625 58.320 129.815 ;
        RECT 58.940 129.675 59.060 129.785 ;
        RECT 59.805 129.645 59.975 129.835 ;
        RECT 62.565 129.625 62.735 129.815 ;
        RECT 64.405 129.625 64.575 129.815 ;
        RECT 65.325 129.645 65.495 129.835 ;
        RECT 69.190 129.645 69.360 129.835 ;
        RECT 71.305 129.645 71.475 129.835 ;
        RECT 73.605 129.815 73.755 129.835 ;
        RECT 73.605 129.645 73.775 129.815 ;
        RECT 74.065 129.625 74.235 129.835 ;
        RECT 74.525 129.645 74.695 129.815 ;
        RECT 76.420 129.675 76.540 129.785 ;
        RECT 76.825 129.645 76.995 129.815 ;
        RECT 78.205 129.645 78.375 129.835 ;
        RECT 80.505 129.815 80.655 129.835 ;
        RECT 80.505 129.645 80.675 129.815 ;
        RECT 74.545 129.625 74.695 129.645 ;
        RECT 76.845 129.625 76.995 129.645 ;
        RECT 82.530 129.625 82.700 129.815 ;
        RECT 83.265 129.645 83.435 129.835 ;
        RECT 85.105 129.645 85.275 129.815 ;
        RECT 85.105 129.625 85.255 129.645 ;
        RECT 86.945 129.625 87.115 129.815 ;
        RECT 87.405 129.625 87.575 129.815 ;
        RECT 88.785 129.645 88.955 129.835 ;
        RECT 89.245 129.785 89.415 129.835 ;
        RECT 89.245 129.675 89.420 129.785 ;
        RECT 89.245 129.645 89.415 129.675 ;
        RECT 89.980 129.625 90.150 129.815 ;
        RECT 93.900 129.675 94.020 129.785 ;
        RECT 94.305 129.625 94.475 129.815 ;
        RECT 95.685 129.625 95.855 129.815 ;
        RECT 101.200 129.645 101.370 129.835 ;
        RECT 102.180 129.675 102.300 129.785 ;
        RECT 103.965 129.645 104.135 129.835 ;
        RECT 106.725 129.645 106.895 129.815 ;
        RECT 109.025 129.645 109.195 129.815 ;
        RECT 109.485 129.645 109.655 129.835 ;
        RECT 111.785 129.815 111.935 129.835 ;
        RECT 111.785 129.645 111.955 129.815 ;
        RECT 112.300 129.675 112.420 129.785 ;
        RECT 113.625 129.645 113.795 129.815 ;
        RECT 115.005 129.785 115.175 129.835 ;
        RECT 114.140 129.675 114.260 129.785 ;
        RECT 115.005 129.675 115.180 129.785 ;
        RECT 115.005 129.645 115.175 129.675 ;
        RECT 106.725 129.625 106.875 129.645 ;
        RECT 109.025 129.625 109.175 129.645 ;
        RECT 14.585 128.815 15.955 129.625 ;
        RECT 15.965 128.815 17.335 129.625 ;
        RECT 17.715 128.945 26.995 129.625 ;
        RECT 17.715 128.825 20.050 128.945 ;
        RECT 17.715 128.715 18.635 128.825 ;
        RECT 24.715 128.725 25.635 128.945 ;
        RECT 27.925 128.815 33.435 129.625 ;
        RECT 33.455 128.715 34.805 129.625 ;
        RECT 35.285 128.815 37.115 129.625 ;
        RECT 37.135 128.755 37.565 129.540 ;
        RECT 38.505 128.845 39.875 129.625 ;
        RECT 40.045 128.805 41.975 129.625 ;
        RECT 42.345 128.805 44.275 129.625 ;
        RECT 45.145 128.815 47.235 129.625 ;
        RECT 47.405 128.805 49.335 129.625 ;
        RECT 49.545 128.815 50.915 129.625 ;
        RECT 50.925 128.815 54.595 129.625 ;
        RECT 54.835 128.945 58.735 129.625 ;
        RECT 41.025 128.715 41.975 128.805 ;
        RECT 43.325 128.715 44.275 128.805 ;
        RECT 48.385 128.715 49.335 128.805 ;
        RECT 57.805 128.715 58.735 128.945 ;
        RECT 59.205 128.815 62.875 129.625 ;
        RECT 62.895 128.755 63.325 129.540 ;
        RECT 63.345 128.815 64.715 129.625 ;
        RECT 65.095 128.945 74.375 129.625 ;
        RECT 65.095 128.825 67.430 128.945 ;
        RECT 65.095 128.715 66.015 128.825 ;
        RECT 72.095 128.725 73.015 128.945 ;
        RECT 74.545 128.805 76.475 129.625 ;
        RECT 76.845 128.805 78.775 129.625 ;
        RECT 79.215 128.945 83.115 129.625 ;
        RECT 75.525 128.715 76.475 128.805 ;
        RECT 77.825 128.715 78.775 128.805 ;
        RECT 82.185 128.715 83.115 128.945 ;
        RECT 83.325 128.805 85.255 129.625 ;
        RECT 85.425 128.815 87.255 129.625 ;
        RECT 87.265 128.845 88.635 129.625 ;
        RECT 83.325 128.715 84.275 128.805 ;
        RECT 88.655 128.755 89.085 129.540 ;
        RECT 89.565 128.945 93.465 129.625 ;
        RECT 89.565 128.715 90.495 128.945 ;
        RECT 94.165 128.845 95.535 129.625 ;
        RECT 95.545 128.945 104.650 129.625 ;
        RECT 104.945 128.805 106.875 129.625 ;
        RECT 107.245 128.805 109.175 129.625 ;
        RECT 109.505 129.625 109.655 129.645 ;
        RECT 113.625 129.625 113.775 129.645 ;
        RECT 117.765 129.625 117.935 129.815 ;
        RECT 118.225 129.625 118.395 129.815 ;
        RECT 119.605 129.625 119.775 129.815 ;
        RECT 120.525 129.645 120.695 129.835 ;
        RECT 126.045 129.625 126.215 129.835 ;
        RECT 127.425 129.625 127.595 129.835 ;
        RECT 109.505 128.805 111.435 129.625 ;
        RECT 104.945 128.715 105.895 128.805 ;
        RECT 107.245 128.715 108.195 128.805 ;
        RECT 110.485 128.715 111.435 128.805 ;
        RECT 111.845 128.805 113.775 129.625 ;
        RECT 111.845 128.715 112.795 128.805 ;
        RECT 114.415 128.755 114.845 129.540 ;
        RECT 115.325 128.815 118.075 129.625 ;
        RECT 118.095 128.715 119.445 129.625 ;
        RECT 119.465 128.845 120.835 129.625 ;
        RECT 120.845 128.815 126.355 129.625 ;
        RECT 126.365 128.815 127.735 129.625 ;
      LAYER nwell ;
        RECT 14.390 125.595 127.930 128.425 ;
      LAYER pwell ;
        RECT 14.585 124.395 15.955 125.205 ;
        RECT 15.965 124.395 17.335 125.205 ;
        RECT 17.345 124.395 21.015 125.205 ;
        RECT 21.035 124.395 22.385 125.305 ;
        RECT 22.865 124.395 24.235 125.175 ;
        RECT 24.255 124.480 24.685 125.265 ;
        RECT 37.805 125.215 38.755 125.305 ;
        RECT 25.625 124.395 31.135 125.205 ;
        RECT 31.145 124.395 36.655 125.205 ;
        RECT 36.825 124.395 38.755 125.215 ;
        RECT 40.545 125.215 41.495 125.305 ;
        RECT 43.785 125.215 44.735 125.305 ;
        RECT 38.965 124.395 40.335 125.205 ;
        RECT 40.545 124.395 42.475 125.215 ;
        RECT 14.725 124.185 14.895 124.395 ;
        RECT 17.025 124.185 17.195 124.395 ;
        RECT 20.705 124.205 20.875 124.395 ;
        RECT 22.085 124.205 22.255 124.395 ;
        RECT 22.545 124.345 22.715 124.375 ;
        RECT 22.545 124.235 22.720 124.345 ;
        RECT 22.545 124.185 22.715 124.235 ;
        RECT 23.005 124.205 23.175 124.395 ;
        RECT 25.305 124.240 25.465 124.350 ;
        RECT 26.410 124.185 26.580 124.375 ;
        RECT 27.200 124.235 27.320 124.345 ;
        RECT 30.825 124.205 30.995 124.395 ;
        RECT 32.665 124.185 32.835 124.375 ;
        RECT 36.345 124.205 36.515 124.395 ;
        RECT 36.825 124.375 36.975 124.395 ;
        RECT 36.530 124.185 36.700 124.375 ;
        RECT 36.805 124.205 36.975 124.375 ;
        RECT 37.780 124.235 37.900 124.345 ;
        RECT 40.025 124.205 40.195 124.395 ;
        RECT 42.325 124.375 42.475 124.395 ;
        RECT 42.805 124.395 44.735 125.215 ;
        RECT 45.145 125.215 46.095 125.305 ;
        RECT 45.145 124.395 47.075 125.215 ;
        RECT 47.255 124.395 49.995 125.075 ;
        RECT 50.015 124.480 50.445 125.265 ;
        RECT 50.465 124.395 52.295 125.205 ;
        RECT 52.305 124.395 57.815 125.205 ;
        RECT 57.825 124.395 59.195 125.175 ;
        RECT 62.405 125.075 63.335 125.305 ;
        RECT 59.435 124.395 63.335 125.075 ;
        RECT 63.345 124.395 64.715 125.205 ;
        RECT 64.725 124.395 68.395 125.205 ;
        RECT 68.415 124.395 69.765 125.305 ;
        RECT 70.245 124.395 71.615 125.175 ;
        RECT 72.545 124.395 75.285 125.075 ;
        RECT 75.775 124.480 76.205 125.265 ;
        RECT 76.225 124.395 78.055 125.205 ;
        RECT 78.435 125.195 79.355 125.305 ;
        RECT 78.435 125.075 80.770 125.195 ;
        RECT 85.435 125.075 86.355 125.295 ;
        RECT 78.435 124.395 87.715 125.075 ;
        RECT 87.725 124.395 89.555 125.205 ;
        RECT 90.925 125.075 91.845 125.295 ;
        RECT 97.925 125.195 98.845 125.305 ;
        RECT 100.365 125.215 101.315 125.305 ;
        RECT 96.510 125.075 98.845 125.195 ;
        RECT 89.565 124.395 98.845 125.075 ;
        RECT 99.385 124.395 101.315 125.215 ;
        RECT 101.535 124.480 101.965 125.265 ;
        RECT 101.985 124.395 105.655 125.205 ;
        RECT 105.665 124.395 111.175 125.205 ;
        RECT 114.385 125.075 115.315 125.305 ;
        RECT 111.415 124.395 115.315 125.075 ;
        RECT 115.695 125.195 116.615 125.305 ;
        RECT 115.695 125.075 118.030 125.195 ;
        RECT 122.695 125.075 123.615 125.295 ;
        RECT 115.695 124.395 124.975 125.075 ;
        RECT 124.985 124.395 126.355 125.205 ;
        RECT 126.365 124.395 127.735 125.205 ;
        RECT 42.805 124.375 42.955 124.395 ;
        RECT 41.405 124.185 41.575 124.375 ;
        RECT 42.325 124.205 42.495 124.375 ;
        RECT 42.785 124.205 42.955 124.375 ;
        RECT 46.925 124.375 47.075 124.395 ;
        RECT 46.925 124.185 47.095 124.375 ;
        RECT 49.685 124.205 49.855 124.395 ;
        RECT 51.985 124.205 52.155 124.395 ;
        RECT 52.445 124.185 52.615 124.375 ;
        RECT 57.505 124.205 57.675 124.395 ;
        RECT 57.965 124.205 58.135 124.395 ;
        RECT 62.105 124.185 62.275 124.375 ;
        RECT 62.620 124.235 62.740 124.345 ;
        RECT 62.750 124.205 62.920 124.395 ;
        RECT 63.540 124.235 63.660 124.345 ;
        RECT 64.405 124.205 64.575 124.395 ;
        RECT 67.350 124.185 67.520 124.375 ;
        RECT 68.085 124.205 68.255 124.395 ;
        RECT 69.465 124.205 69.635 124.395 ;
        RECT 69.980 124.235 70.100 124.345 ;
        RECT 70.385 124.185 70.555 124.395 ;
        RECT 72.225 124.240 72.385 124.350 ;
        RECT 72.685 124.205 72.855 124.395 ;
        RECT 75.500 124.235 75.620 124.345 ;
        RECT 75.905 124.185 76.075 124.375 ;
        RECT 77.745 124.205 77.915 124.395 ;
        RECT 81.425 124.185 81.595 124.375 ;
        RECT 82.805 124.185 82.975 124.375 ;
        RECT 83.320 124.235 83.440 124.345 ;
        RECT 83.725 124.185 83.895 124.375 ;
        RECT 87.405 124.205 87.575 124.395 ;
        RECT 88.325 124.185 88.495 124.375 ;
        RECT 89.245 124.205 89.415 124.395 ;
        RECT 89.705 124.205 89.875 124.395 ;
        RECT 99.385 124.375 99.535 124.395 ;
        RECT 92.465 124.185 92.635 124.375 ;
        RECT 92.925 124.185 93.095 124.375 ;
        RECT 95.225 124.185 95.395 124.375 ;
        RECT 98.905 124.185 99.075 124.375 ;
        RECT 99.365 124.205 99.535 124.375 ;
        RECT 104.425 124.185 104.595 124.375 ;
        RECT 105.345 124.205 105.515 124.395 ;
        RECT 109.945 124.185 110.115 124.375 ;
        RECT 110.865 124.205 111.035 124.395 ;
        RECT 113.810 124.185 113.980 124.375 ;
        RECT 114.730 124.205 114.900 124.395 ;
        RECT 115.060 124.235 115.180 124.345 ;
        RECT 124.665 124.185 124.835 124.395 ;
        RECT 126.045 124.185 126.215 124.395 ;
        RECT 127.425 124.185 127.595 124.395 ;
        RECT 14.585 123.375 15.955 124.185 ;
        RECT 15.965 123.375 17.335 124.185 ;
        RECT 17.345 123.375 22.855 124.185 ;
        RECT 23.095 123.505 26.995 124.185 ;
        RECT 26.065 123.275 26.995 123.505 ;
        RECT 27.465 123.375 32.975 124.185 ;
        RECT 33.215 123.505 37.115 124.185 ;
        RECT 36.185 123.275 37.115 123.505 ;
        RECT 37.135 123.315 37.565 124.100 ;
        RECT 38.045 123.375 41.715 124.185 ;
        RECT 41.725 123.375 47.235 124.185 ;
        RECT 47.245 123.375 52.755 124.185 ;
        RECT 53.135 123.505 62.415 124.185 ;
        RECT 53.135 123.385 55.470 123.505 ;
        RECT 53.135 123.275 54.055 123.385 ;
        RECT 60.135 123.285 61.055 123.505 ;
        RECT 62.895 123.315 63.325 124.100 ;
        RECT 64.035 123.505 67.935 124.185 ;
        RECT 67.005 123.275 67.935 123.505 ;
        RECT 67.945 123.375 70.695 124.185 ;
        RECT 70.705 123.375 76.215 124.185 ;
        RECT 76.225 123.375 81.735 124.185 ;
        RECT 81.755 123.275 83.105 124.185 ;
        RECT 83.585 123.405 84.955 124.185 ;
        RECT 84.965 123.375 88.635 124.185 ;
        RECT 88.655 123.315 89.085 124.100 ;
        RECT 89.105 123.375 92.775 124.185 ;
        RECT 92.795 123.275 94.145 124.185 ;
        RECT 94.165 123.375 95.535 124.185 ;
        RECT 95.545 123.375 99.215 124.185 ;
        RECT 99.225 123.375 104.735 124.185 ;
        RECT 104.745 123.375 110.255 124.185 ;
        RECT 110.495 123.505 114.395 124.185 ;
        RECT 113.465 123.275 114.395 123.505 ;
        RECT 114.415 123.315 114.845 124.100 ;
        RECT 115.695 123.505 124.975 124.185 ;
        RECT 115.695 123.385 118.030 123.505 ;
        RECT 115.695 123.275 116.615 123.385 ;
        RECT 122.695 123.285 123.615 123.505 ;
        RECT 124.985 123.375 126.355 124.185 ;
        RECT 126.365 123.375 127.735 124.185 ;
      LAYER nwell ;
        RECT 14.390 120.155 127.930 122.985 ;
      LAYER pwell ;
        RECT 14.585 118.955 15.955 119.765 ;
        RECT 16.425 118.955 20.095 119.765 ;
        RECT 20.105 119.635 21.035 119.865 ;
        RECT 20.105 118.955 24.005 119.635 ;
        RECT 24.255 119.040 24.685 119.825 ;
        RECT 24.705 118.955 26.075 119.765 ;
        RECT 26.085 118.955 27.455 119.735 ;
        RECT 27.465 118.955 30.215 119.765 ;
        RECT 30.595 119.755 31.515 119.865 ;
        RECT 30.595 119.635 32.930 119.755 ;
        RECT 37.595 119.635 38.515 119.855 ;
        RECT 39.885 119.635 40.815 119.865 ;
        RECT 30.595 118.955 39.875 119.635 ;
        RECT 39.885 118.955 43.785 119.635 ;
        RECT 44.485 118.955 45.855 119.735 ;
        RECT 49.065 119.635 49.995 119.865 ;
        RECT 46.095 118.955 49.995 119.635 ;
        RECT 50.015 119.040 50.445 119.825 ;
        RECT 50.475 118.955 51.825 119.865 ;
        RECT 51.845 118.955 53.215 119.765 ;
        RECT 53.365 118.955 55.975 119.865 ;
        RECT 56.915 118.955 58.265 119.865 ;
        RECT 59.575 119.755 60.495 119.865 ;
        RECT 59.575 119.635 61.910 119.755 ;
        RECT 66.575 119.635 67.495 119.855 ;
        RECT 59.575 118.955 68.855 119.635 ;
        RECT 68.865 118.955 70.235 119.735 ;
        RECT 70.705 118.955 74.375 119.765 ;
        RECT 74.395 118.955 75.745 119.865 ;
        RECT 75.775 119.040 76.205 119.825 ;
        RECT 79.885 119.635 80.815 119.865 ;
        RECT 76.915 118.955 80.815 119.635 ;
        RECT 80.825 118.955 82.195 119.735 ;
        RECT 82.215 118.955 83.565 119.865 ;
        RECT 84.045 118.955 85.415 119.735 ;
        RECT 85.425 118.955 90.935 119.765 ;
        RECT 90.945 119.635 91.875 119.865 ;
        RECT 90.945 118.955 94.845 119.635 ;
        RECT 95.545 118.955 97.375 119.765 ;
        RECT 100.585 119.635 101.515 119.865 ;
        RECT 97.615 118.955 101.515 119.635 ;
        RECT 101.535 119.040 101.965 119.825 ;
        RECT 101.985 118.955 103.355 119.765 ;
        RECT 103.375 118.955 104.725 119.865 ;
        RECT 107.945 119.635 108.875 119.865 ;
        RECT 104.975 118.955 108.875 119.635 ;
        RECT 109.255 119.755 110.175 119.865 ;
        RECT 109.255 119.635 111.590 119.755 ;
        RECT 116.255 119.635 117.175 119.855 ;
        RECT 109.255 118.955 118.535 119.635 ;
        RECT 118.555 118.955 119.905 119.865 ;
        RECT 120.385 118.955 121.755 119.735 ;
        RECT 122.685 118.955 126.355 119.765 ;
        RECT 126.365 118.955 127.735 119.765 ;
        RECT 14.725 118.745 14.895 118.955 ;
        RECT 16.160 118.795 16.280 118.905 ;
        RECT 17.485 118.745 17.655 118.935 ;
        RECT 19.785 118.765 19.955 118.955 ;
        RECT 20.520 118.765 20.690 118.955 ;
        RECT 25.765 118.765 25.935 118.955 ;
        RECT 27.145 118.745 27.315 118.955 ;
        RECT 27.605 118.745 27.775 118.935 ;
        RECT 29.905 118.765 30.075 118.955 ;
        RECT 39.565 118.765 39.735 118.955 ;
        RECT 40.300 118.765 40.470 118.955 ;
        RECT 44.220 118.795 44.340 118.905 ;
        RECT 45.545 118.765 45.715 118.955 ;
        RECT 46.925 118.745 47.095 118.935 ;
        RECT 49.410 118.765 49.580 118.955 ;
        RECT 50.605 118.765 50.775 118.955 ;
        RECT 52.905 118.765 53.075 118.955 ;
        RECT 55.660 118.765 55.830 118.955 ;
        RECT 56.585 118.745 56.755 118.935 ;
        RECT 57.505 118.790 57.665 118.900 ;
        RECT 57.965 118.765 58.135 118.955 ;
        RECT 58.885 118.800 59.045 118.910 ;
        RECT 61.185 118.745 61.355 118.935 ;
        RECT 61.645 118.745 61.815 118.935 ;
        RECT 68.545 118.765 68.715 118.955 ;
        RECT 69.925 118.765 70.095 118.955 ;
        RECT 70.440 118.795 70.560 118.905 ;
        RECT 72.685 118.745 72.855 118.935 ;
        RECT 74.065 118.765 74.235 118.955 ;
        RECT 74.525 118.765 74.695 118.955 ;
        RECT 76.420 118.795 76.540 118.905 ;
        RECT 80.230 118.765 80.400 118.955 ;
        RECT 81.885 118.765 82.055 118.955 ;
        RECT 82.345 118.745 82.515 118.935 ;
        RECT 83.080 118.745 83.250 118.935 ;
        RECT 83.265 118.765 83.435 118.955 ;
        RECT 83.780 118.795 83.900 118.905 ;
        RECT 84.185 118.765 84.355 118.955 ;
        RECT 87.000 118.795 87.120 118.905 ;
        RECT 87.405 118.745 87.575 118.935 ;
        RECT 89.245 118.745 89.415 118.935 ;
        RECT 90.625 118.745 90.795 118.955 ;
        RECT 91.360 118.765 91.530 118.955 ;
        RECT 92.465 118.790 92.625 118.900 ;
        RECT 95.280 118.795 95.400 118.905 ;
        RECT 97.065 118.765 97.235 118.955 ;
        RECT 100.930 118.765 101.100 118.955 ;
        RECT 102.125 118.745 102.295 118.935 ;
        RECT 103.045 118.765 103.215 118.955 ;
        RECT 103.505 118.765 103.675 118.955 ;
        RECT 108.290 118.765 108.460 118.955 ;
        RECT 111.785 118.745 111.955 118.935 ;
        RECT 112.705 118.790 112.865 118.900 ;
        RECT 114.085 118.745 114.255 118.935 ;
        RECT 115.060 118.795 115.180 118.905 ;
        RECT 115.465 118.745 115.635 118.935 ;
        RECT 116.900 118.795 117.020 118.905 ;
        RECT 118.225 118.765 118.395 118.955 ;
        RECT 118.685 118.765 118.855 118.955 ;
        RECT 120.120 118.795 120.240 118.905 ;
        RECT 120.525 118.745 120.695 118.955 ;
        RECT 122.365 118.800 122.525 118.910 ;
        RECT 126.045 118.745 126.215 118.955 ;
        RECT 127.425 118.745 127.595 118.955 ;
        RECT 14.585 117.935 15.955 118.745 ;
        RECT 16.435 117.835 17.785 118.745 ;
        RECT 18.175 118.065 27.455 118.745 ;
        RECT 27.465 118.065 36.745 118.745 ;
        RECT 18.175 117.945 20.510 118.065 ;
        RECT 18.175 117.835 19.095 117.945 ;
        RECT 25.175 117.845 26.095 118.065 ;
        RECT 28.825 117.845 29.745 118.065 ;
        RECT 34.410 117.945 36.745 118.065 ;
        RECT 35.825 117.835 36.745 117.945 ;
        RECT 37.135 117.875 37.565 118.660 ;
        RECT 37.955 118.065 47.235 118.745 ;
        RECT 47.615 118.065 56.895 118.745 ;
        RECT 37.955 117.945 40.290 118.065 ;
        RECT 37.955 117.835 38.875 117.945 ;
        RECT 44.955 117.845 45.875 118.065 ;
        RECT 47.615 117.945 49.950 118.065 ;
        RECT 47.615 117.835 48.535 117.945 ;
        RECT 54.615 117.845 55.535 118.065 ;
        RECT 57.825 117.935 61.495 118.745 ;
        RECT 61.515 117.835 62.865 118.745 ;
        RECT 62.895 117.875 63.325 118.660 ;
        RECT 63.715 118.065 72.995 118.745 ;
        RECT 73.375 118.065 82.655 118.745 ;
        RECT 82.665 118.065 86.565 118.745 ;
        RECT 63.715 117.945 66.050 118.065 ;
        RECT 63.715 117.835 64.635 117.945 ;
        RECT 70.715 117.845 71.635 118.065 ;
        RECT 73.375 117.945 75.710 118.065 ;
        RECT 73.375 117.835 74.295 117.945 ;
        RECT 80.375 117.845 81.295 118.065 ;
        RECT 82.665 117.835 83.595 118.065 ;
        RECT 87.265 117.965 88.635 118.745 ;
        RECT 88.655 117.875 89.085 118.660 ;
        RECT 89.115 117.835 90.465 118.745 ;
        RECT 90.495 117.835 91.845 118.745 ;
        RECT 93.155 118.065 102.435 118.745 ;
        RECT 102.815 118.065 112.095 118.745 ;
        RECT 93.155 117.945 95.490 118.065 ;
        RECT 93.155 117.835 94.075 117.945 ;
        RECT 100.155 117.845 101.075 118.065 ;
        RECT 102.815 117.945 105.150 118.065 ;
        RECT 102.815 117.835 103.735 117.945 ;
        RECT 109.815 117.845 110.735 118.065 ;
        RECT 113.035 117.835 114.385 118.745 ;
        RECT 114.415 117.875 114.845 118.660 ;
        RECT 115.325 117.965 116.695 118.745 ;
        RECT 117.165 117.935 120.835 118.745 ;
        RECT 120.845 117.935 126.355 118.745 ;
        RECT 126.365 117.935 127.735 118.745 ;
      LAYER nwell ;
        RECT 14.390 114.715 127.930 117.545 ;
      LAYER pwell ;
        RECT 14.585 113.515 15.955 114.325 ;
        RECT 15.965 113.515 17.335 114.325 ;
        RECT 17.345 113.515 21.015 114.325 ;
        RECT 21.025 113.515 22.395 114.295 ;
        RECT 22.415 113.515 23.765 114.425 ;
        RECT 24.255 113.600 24.685 114.385 ;
        RECT 26.065 114.195 26.985 114.415 ;
        RECT 33.065 114.315 33.985 114.425 ;
        RECT 31.650 114.195 33.985 114.315 ;
        RECT 24.705 113.515 33.985 114.195 ;
        RECT 34.835 113.515 36.185 114.425 ;
        RECT 36.665 113.515 38.035 114.295 ;
        RECT 38.965 113.515 40.335 114.295 ;
        RECT 40.345 113.515 44.015 114.325 ;
        RECT 44.035 113.515 45.385 114.425 ;
        RECT 45.405 114.195 46.335 114.425 ;
        RECT 45.405 113.515 49.305 114.195 ;
        RECT 50.015 113.600 50.445 114.385 ;
        RECT 50.465 113.515 52.295 114.325 ;
        RECT 52.305 113.515 53.675 114.295 ;
        RECT 53.685 113.515 55.055 114.325 ;
        RECT 55.065 113.515 60.575 114.325 ;
        RECT 60.585 113.515 66.095 114.325 ;
        RECT 66.115 113.515 67.465 114.425 ;
        RECT 67.945 113.515 69.315 114.295 ;
        RECT 70.245 113.515 75.755 114.325 ;
        RECT 75.775 113.600 76.205 114.385 ;
        RECT 77.515 114.315 78.435 114.425 ;
        RECT 77.515 114.195 79.850 114.315 ;
        RECT 84.515 114.195 85.435 114.415 ;
        RECT 88.625 114.195 89.545 114.415 ;
        RECT 95.625 114.315 96.545 114.425 ;
        RECT 94.210 114.195 96.545 114.315 ;
        RECT 77.515 113.515 86.795 114.195 ;
        RECT 87.265 113.515 96.545 114.195 ;
        RECT 97.385 113.515 100.135 114.325 ;
        RECT 100.145 113.515 101.515 114.295 ;
        RECT 101.535 113.600 101.965 114.385 ;
        RECT 102.445 113.515 107.955 114.325 ;
        RECT 107.965 113.515 109.335 114.295 ;
        RECT 109.345 113.515 111.175 114.325 ;
        RECT 114.385 114.195 115.315 114.425 ;
        RECT 111.415 113.515 115.315 114.195 ;
        RECT 115.325 113.515 120.835 114.325 ;
        RECT 120.845 113.515 126.355 114.325 ;
        RECT 126.365 113.515 127.735 114.325 ;
        RECT 14.725 113.305 14.895 113.515 ;
        RECT 17.025 113.325 17.195 113.515 ;
        RECT 20.705 113.325 20.875 113.515 ;
        RECT 21.165 113.325 21.335 113.515 ;
        RECT 23.465 113.325 23.635 113.515 ;
        RECT 23.980 113.355 24.100 113.465 ;
        RECT 24.845 113.325 25.015 113.515 ;
        RECT 26.225 113.305 26.395 113.495 ;
        RECT 28.065 113.305 28.235 113.495 ;
        RECT 33.585 113.305 33.755 113.495 ;
        RECT 34.560 113.355 34.680 113.465 ;
        RECT 34.965 113.305 35.135 113.495 ;
        RECT 35.885 113.325 36.055 113.515 ;
        RECT 36.400 113.355 36.520 113.465 ;
        RECT 36.805 113.305 36.975 113.515 ;
        RECT 37.780 113.355 37.900 113.465 ;
        RECT 38.645 113.360 38.805 113.470 ;
        RECT 40.025 113.325 40.195 113.515 ;
        RECT 43.705 113.325 43.875 113.515 ;
        RECT 45.085 113.325 45.255 113.515 ;
        RECT 45.820 113.325 45.990 113.515 ;
        RECT 46.925 113.305 47.095 113.495 ;
        RECT 47.845 113.350 48.005 113.460 ;
        RECT 49.740 113.355 49.860 113.465 ;
        RECT 51.525 113.305 51.695 113.495 ;
        RECT 51.985 113.325 52.155 113.515 ;
        RECT 52.445 113.325 52.615 113.515 ;
        RECT 54.745 113.325 54.915 113.515 ;
        RECT 57.045 113.305 57.215 113.495 ;
        RECT 60.265 113.325 60.435 113.515 ;
        RECT 62.565 113.305 62.735 113.495 ;
        RECT 63.540 113.355 63.660 113.465 ;
        RECT 65.785 113.325 65.955 113.515 ;
        RECT 66.245 113.325 66.415 113.515 ;
        RECT 67.680 113.355 67.800 113.465 ;
        RECT 68.085 113.325 68.255 113.515 ;
        RECT 69.005 113.305 69.175 113.495 ;
        RECT 69.925 113.360 70.085 113.470 ;
        RECT 74.525 113.305 74.695 113.495 ;
        RECT 75.445 113.325 75.615 113.515 ;
        RECT 76.825 113.360 76.985 113.470 ;
        RECT 80.045 113.305 80.215 113.495 ;
        RECT 81.425 113.305 81.595 113.495 ;
        RECT 82.805 113.305 82.975 113.495 ;
        RECT 86.485 113.325 86.655 113.515 ;
        RECT 87.000 113.355 87.120 113.465 ;
        RECT 87.405 113.325 87.575 113.515 ;
        RECT 88.325 113.305 88.495 113.495 ;
        RECT 92.465 113.305 92.635 113.495 ;
        RECT 92.925 113.305 93.095 113.495 ;
        RECT 97.120 113.355 97.240 113.465 ;
        RECT 99.825 113.325 99.995 113.515 ;
        RECT 101.205 113.325 101.375 113.515 ;
        RECT 102.180 113.355 102.300 113.465 ;
        RECT 103.045 113.325 103.215 113.495 ;
        RECT 107.645 113.325 107.815 113.515 ;
        RECT 108.105 113.325 108.275 113.515 ;
        RECT 108.565 113.305 108.735 113.495 ;
        RECT 110.865 113.325 111.035 113.515 ;
        RECT 114.085 113.305 114.255 113.495 ;
        RECT 114.730 113.325 114.900 113.515 ;
        RECT 115.465 113.350 115.625 113.460 ;
        RECT 119.145 113.305 119.315 113.495 ;
        RECT 119.605 113.305 119.775 113.495 ;
        RECT 120.525 113.325 120.695 113.515 ;
        RECT 121.905 113.305 122.075 113.495 ;
        RECT 123.285 113.305 123.455 113.495 ;
        RECT 126.045 113.305 126.215 113.515 ;
        RECT 127.425 113.305 127.595 113.515 ;
        RECT 14.585 112.495 15.955 113.305 ;
        RECT 16.165 112.625 26.535 113.305 ;
        RECT 16.165 112.395 18.375 112.625 ;
        RECT 21.095 112.405 22.025 112.625 ;
        RECT 26.545 112.495 28.375 113.305 ;
        RECT 28.385 112.495 33.895 113.305 ;
        RECT 33.915 112.395 35.265 113.305 ;
        RECT 35.285 112.495 37.115 113.305 ;
        RECT 37.135 112.435 37.565 113.220 ;
        RECT 38.130 112.625 47.235 113.305 ;
        RECT 48.165 112.495 51.835 113.305 ;
        RECT 51.845 112.495 57.355 113.305 ;
        RECT 57.365 112.495 62.875 113.305 ;
        RECT 62.895 112.435 63.325 113.220 ;
        RECT 63.805 112.495 69.315 113.305 ;
        RECT 69.325 112.495 74.835 113.305 ;
        RECT 74.845 112.495 80.355 113.305 ;
        RECT 80.375 112.395 81.725 113.305 ;
        RECT 81.745 112.495 83.115 113.305 ;
        RECT 83.125 112.495 88.635 113.305 ;
        RECT 88.655 112.435 89.085 113.220 ;
        RECT 89.105 112.495 92.775 113.305 ;
        RECT 92.785 112.625 101.890 113.305 ;
        RECT 101.985 112.625 102.940 113.305 ;
        RECT 103.365 112.495 108.875 113.305 ;
        RECT 108.885 112.495 114.395 113.305 ;
        RECT 114.415 112.435 114.845 113.220 ;
        RECT 115.785 112.495 119.455 113.305 ;
        RECT 119.475 112.395 120.825 113.305 ;
        RECT 120.845 112.525 122.215 113.305 ;
        RECT 122.225 112.525 123.595 113.305 ;
        RECT 123.605 112.495 126.355 113.305 ;
        RECT 126.365 112.495 127.735 113.305 ;
      LAYER nwell ;
        RECT 14.390 109.275 127.930 112.105 ;
      LAYER pwell ;
        RECT 14.585 108.075 15.955 108.885 ;
        RECT 16.885 108.075 20.555 108.885 ;
        RECT 20.575 108.075 21.925 108.985 ;
        RECT 22.875 108.075 24.225 108.985 ;
        RECT 24.255 108.160 24.685 108.945 ;
        RECT 24.705 108.075 27.455 108.885 ;
        RECT 27.465 108.075 28.835 108.855 ;
        RECT 28.845 108.075 30.675 108.885 ;
        RECT 30.695 108.075 32.045 108.985 ;
        RECT 32.065 108.075 33.435 108.855 ;
        RECT 34.365 108.075 35.735 108.855 ;
        RECT 36.205 108.075 38.955 108.885 ;
        RECT 38.965 108.075 44.475 108.885 ;
        RECT 44.485 108.075 49.995 108.885 ;
        RECT 50.015 108.160 50.445 108.945 ;
        RECT 50.925 108.075 52.295 108.855 ;
        RECT 53.225 108.075 56.895 108.885 ;
        RECT 56.905 108.075 58.275 108.855 ;
        RECT 58.285 108.075 59.655 108.885 ;
        RECT 59.665 108.075 62.275 108.985 ;
        RECT 62.885 108.075 64.715 108.885 ;
        RECT 64.735 108.075 66.085 108.985 ;
        RECT 66.565 108.075 68.395 108.885 ;
        RECT 68.405 108.075 69.775 108.855 ;
        RECT 70.245 108.075 75.755 108.885 ;
        RECT 75.775 108.160 76.205 108.945 ;
        RECT 76.235 108.075 77.585 108.985 ;
        RECT 77.615 108.075 78.965 108.985 ;
        RECT 79.905 108.075 82.515 108.985 ;
        RECT 82.665 108.075 84.035 108.855 ;
        RECT 84.505 108.075 87.255 108.885 ;
        RECT 87.275 108.075 88.625 108.985 ;
        RECT 88.645 108.075 92.315 108.885 ;
        RECT 92.335 108.075 93.685 108.985 ;
        RECT 93.705 108.075 95.075 108.855 ;
        RECT 95.085 108.075 96.455 108.885 ;
        RECT 96.465 108.075 100.135 108.885 ;
        RECT 100.145 108.075 101.515 108.855 ;
        RECT 101.535 108.160 101.965 108.945 ;
        RECT 102.445 108.075 106.115 108.885 ;
        RECT 106.125 108.075 107.495 108.855 ;
        RECT 107.505 108.075 108.875 108.885 ;
        RECT 108.895 108.075 110.245 108.985 ;
        RECT 110.265 108.075 111.635 108.855 ;
        RECT 111.645 108.075 113.015 108.855 ;
        RECT 113.025 108.075 114.395 108.885 ;
        RECT 114.415 108.075 115.765 108.985 ;
        RECT 120.295 108.755 121.225 108.975 ;
        RECT 123.945 108.755 126.155 108.985 ;
        RECT 115.785 108.075 126.155 108.755 ;
        RECT 126.365 108.075 127.735 108.885 ;
        RECT 14.725 107.865 14.895 108.075 ;
        RECT 16.565 107.920 16.725 108.030 ;
        RECT 20.245 107.885 20.415 108.075 ;
        RECT 21.625 107.885 21.795 108.075 ;
        RECT 22.545 107.920 22.705 108.030 ;
        RECT 23.925 107.885 24.095 108.075 ;
        RECT 26.225 107.865 26.395 108.055 ;
        RECT 27.145 107.885 27.315 108.075 ;
        RECT 28.525 107.885 28.695 108.075 ;
        RECT 30.365 107.885 30.535 108.075 ;
        RECT 31.745 107.885 31.915 108.075 ;
        RECT 33.125 107.885 33.295 108.075 ;
        RECT 34.045 107.920 34.205 108.030 ;
        RECT 35.425 107.885 35.595 108.075 ;
        RECT 35.940 107.915 36.060 108.025 ;
        RECT 36.805 107.865 36.975 108.055 ;
        RECT 38.645 107.865 38.815 108.075 ;
        RECT 39.160 107.915 39.280 108.025 ;
        RECT 40.485 107.865 40.655 108.055 ;
        RECT 41.865 107.865 42.035 108.055 ;
        RECT 43.245 107.865 43.415 108.055 ;
        RECT 43.760 107.915 43.880 108.025 ;
        RECT 44.165 107.885 44.335 108.075 ;
        RECT 45.085 107.865 45.255 108.055 ;
        RECT 45.545 107.865 45.715 108.055 ;
        RECT 49.685 107.885 49.855 108.075 ;
        RECT 50.660 107.915 50.780 108.025 ;
        RECT 51.065 107.885 51.235 108.075 ;
        RECT 52.905 107.920 53.065 108.030 ;
        RECT 56.585 107.885 56.755 108.075 ;
        RECT 57.045 107.865 57.215 108.075 ;
        RECT 58.425 107.865 58.595 108.055 ;
        RECT 59.345 107.885 59.515 108.075 ;
        RECT 59.810 108.055 59.980 108.075 ;
        RECT 59.805 107.885 59.980 108.055 ;
        RECT 59.805 107.865 59.975 107.885 ;
        RECT 60.265 107.865 60.435 108.055 ;
        RECT 61.645 107.865 61.815 108.055 ;
        RECT 62.620 107.915 62.740 108.025 ;
        RECT 64.405 107.885 64.575 108.075 ;
        RECT 64.865 107.885 65.035 108.075 ;
        RECT 66.300 107.915 66.420 108.025 ;
        RECT 68.085 107.885 68.255 108.075 ;
        RECT 68.545 107.885 68.715 108.075 ;
        RECT 69.980 107.915 70.100 108.025 ;
        RECT 73.605 107.865 73.775 108.055 ;
        RECT 74.525 107.910 74.685 108.020 ;
        RECT 74.985 107.865 75.155 108.055 ;
        RECT 75.445 107.885 75.615 108.075 ;
        RECT 77.285 107.885 77.455 108.075 ;
        RECT 78.665 107.885 78.835 108.075 ;
        RECT 79.585 107.920 79.745 108.030 ;
        RECT 80.050 107.885 80.220 108.075 ;
        RECT 82.805 107.885 82.975 108.075 ;
        RECT 84.240 107.915 84.360 108.025 ;
        RECT 86.485 107.865 86.655 108.055 ;
        RECT 86.945 108.025 87.115 108.075 ;
        RECT 86.945 107.915 87.120 108.025 ;
        RECT 86.945 107.885 87.115 107.915 ;
        RECT 87.405 107.865 87.575 108.075 ;
        RECT 92.005 107.885 92.175 108.075 ;
        RECT 92.465 107.885 92.635 108.075 ;
        RECT 93.845 107.885 94.015 108.075 ;
        RECT 96.145 107.885 96.315 108.075 ;
        RECT 99.365 107.865 99.535 108.055 ;
        RECT 99.825 107.885 99.995 108.075 ;
        RECT 100.745 107.865 100.915 108.055 ;
        RECT 101.205 107.885 101.375 108.075 ;
        RECT 102.125 108.025 102.295 108.055 ;
        RECT 102.125 107.915 102.300 108.025 ;
        RECT 102.125 107.865 102.295 107.915 ;
        RECT 102.585 107.865 102.755 108.055 ;
        RECT 105.805 107.885 105.975 108.075 ;
        RECT 106.265 107.885 106.435 108.075 ;
        RECT 108.565 107.885 108.735 108.075 ;
        RECT 109.945 107.885 110.115 108.075 ;
        RECT 110.405 107.885 110.575 108.075 ;
        RECT 111.785 107.885 111.955 108.075 ;
        RECT 114.085 107.865 114.255 108.075 ;
        RECT 114.545 107.885 114.715 108.075 ;
        RECT 115.465 107.910 115.625 108.020 ;
        RECT 115.925 107.865 116.095 108.075 ;
        RECT 127.425 107.865 127.595 108.075 ;
        RECT 14.585 107.055 15.955 107.865 ;
        RECT 16.165 107.185 26.535 107.865 ;
        RECT 26.745 107.185 37.115 107.865 ;
        RECT 16.165 106.955 18.375 107.185 ;
        RECT 21.095 106.965 22.025 107.185 ;
        RECT 26.745 106.955 28.955 107.185 ;
        RECT 31.675 106.965 32.605 107.185 ;
        RECT 37.135 106.995 37.565 107.780 ;
        RECT 37.585 107.085 38.955 107.865 ;
        RECT 39.435 106.955 40.785 107.865 ;
        RECT 40.805 107.055 42.175 107.865 ;
        RECT 42.185 107.085 43.555 107.865 ;
        RECT 44.035 106.955 45.385 107.865 ;
        RECT 45.405 107.085 46.775 107.865 ;
        RECT 46.985 107.185 57.355 107.865 ;
        RECT 46.985 106.955 49.195 107.185 ;
        RECT 51.915 106.965 52.845 107.185 ;
        RECT 57.375 106.955 58.725 107.865 ;
        RECT 58.745 107.055 60.115 107.865 ;
        RECT 60.135 106.955 61.485 107.865 ;
        RECT 61.505 107.085 62.875 107.865 ;
        RECT 62.895 106.995 63.325 107.780 ;
        RECT 63.545 107.185 73.915 107.865 ;
        RECT 63.545 106.955 65.755 107.185 ;
        RECT 68.475 106.965 69.405 107.185 ;
        RECT 74.845 107.085 76.215 107.865 ;
        RECT 76.425 107.185 86.795 107.865 ;
        RECT 76.425 106.955 78.635 107.185 ;
        RECT 81.355 106.965 82.285 107.185 ;
        RECT 87.265 107.085 88.635 107.865 ;
        RECT 88.655 106.995 89.085 107.780 ;
        RECT 89.305 107.185 99.675 107.865 ;
        RECT 89.305 106.955 91.515 107.185 ;
        RECT 94.235 106.965 95.165 107.185 ;
        RECT 99.695 106.955 101.045 107.865 ;
        RECT 101.065 107.055 102.435 107.865 ;
        RECT 102.455 106.955 103.805 107.865 ;
        RECT 104.025 107.185 114.395 107.865 ;
        RECT 104.025 106.955 106.235 107.185 ;
        RECT 108.955 106.965 109.885 107.185 ;
        RECT 114.415 106.995 114.845 107.780 ;
        RECT 115.785 107.185 126.155 107.865 ;
        RECT 120.295 106.965 121.225 107.185 ;
        RECT 123.945 106.955 126.155 107.185 ;
        RECT 126.365 107.055 127.735 107.865 ;
      LAYER nwell ;
        RECT 14.390 103.835 127.930 106.665 ;
      LAYER pwell ;
        RECT 14.585 102.635 15.955 103.445 ;
        RECT 15.965 102.635 18.715 103.445 ;
        RECT 18.725 102.635 24.235 103.445 ;
        RECT 24.255 102.720 24.685 103.505 ;
        RECT 24.705 102.635 27.455 103.445 ;
        RECT 27.475 102.635 28.825 103.545 ;
        RECT 33.355 103.315 34.285 103.535 ;
        RECT 37.005 103.315 39.215 103.545 ;
        RECT 28.845 102.635 39.215 103.315 ;
        RECT 39.625 103.315 41.835 103.545 ;
        RECT 44.555 103.315 45.485 103.535 ;
        RECT 39.625 102.635 49.995 103.315 ;
        RECT 50.015 102.720 50.445 103.505 ;
        RECT 51.395 102.635 52.745 103.545 ;
        RECT 52.965 103.315 55.175 103.545 ;
        RECT 57.895 103.315 58.825 103.535 ;
        RECT 63.545 103.315 65.755 103.545 ;
        RECT 68.475 103.315 69.405 103.535 ;
        RECT 52.965 102.635 63.335 103.315 ;
        RECT 63.545 102.635 73.915 103.315 ;
        RECT 73.925 102.635 75.755 103.445 ;
        RECT 75.775 102.720 76.205 103.505 ;
        RECT 76.425 103.315 78.635 103.545 ;
        RECT 81.355 103.315 82.285 103.535 ;
        RECT 87.005 103.315 89.215 103.545 ;
        RECT 91.935 103.315 92.865 103.535 ;
        RECT 76.425 102.635 86.795 103.315 ;
        RECT 87.005 102.635 97.375 103.315 ;
        RECT 97.845 102.635 101.515 103.445 ;
        RECT 101.535 102.720 101.965 103.505 ;
        RECT 102.185 103.315 104.395 103.545 ;
        RECT 107.115 103.315 108.045 103.535 ;
        RECT 117.075 103.315 118.005 103.535 ;
        RECT 120.725 103.315 122.935 103.545 ;
        RECT 102.185 102.635 112.555 103.315 ;
        RECT 112.565 102.635 122.935 103.315 ;
        RECT 123.145 102.635 124.975 103.445 ;
        RECT 124.985 102.635 126.355 103.415 ;
        RECT 126.365 102.635 127.735 103.445 ;
        RECT 14.725 102.425 14.895 102.635 ;
        RECT 18.405 102.425 18.575 102.635 ;
        RECT 23.925 102.425 24.095 102.635 ;
        RECT 27.145 102.445 27.315 102.635 ;
        RECT 27.605 102.445 27.775 102.635 ;
        RECT 28.985 102.445 29.155 102.635 ;
        RECT 34.965 102.425 35.135 102.615 ;
        RECT 36.805 102.425 36.975 102.615 ;
        RECT 38.645 102.425 38.815 102.615 ;
        RECT 44.165 102.425 44.335 102.615 ;
        RECT 49.685 102.425 49.855 102.635 ;
        RECT 51.065 102.480 51.225 102.590 ;
        RECT 51.525 102.425 51.695 102.615 ;
        RECT 52.445 102.445 52.615 102.635 ;
        RECT 57.045 102.425 57.215 102.615 ;
        RECT 62.565 102.425 62.735 102.615 ;
        RECT 63.025 102.445 63.195 102.635 ;
        RECT 64.405 102.425 64.575 102.615 ;
        RECT 69.925 102.425 70.095 102.615 ;
        RECT 73.605 102.445 73.775 102.635 ;
        RECT 75.445 102.425 75.615 102.635 ;
        RECT 77.285 102.425 77.455 102.615 ;
        RECT 82.805 102.425 82.975 102.615 ;
        RECT 86.485 102.445 86.655 102.635 ;
        RECT 88.325 102.425 88.495 102.615 ;
        RECT 90.625 102.425 90.795 102.615 ;
        RECT 97.065 102.445 97.235 102.635 ;
        RECT 97.580 102.475 97.700 102.585 ;
        RECT 101.205 102.425 101.375 102.635 ;
        RECT 103.045 102.425 103.215 102.615 ;
        RECT 108.565 102.425 108.735 102.615 ;
        RECT 112.245 102.445 112.415 102.635 ;
        RECT 112.705 102.445 112.875 102.635 ;
        RECT 114.085 102.425 114.255 102.615 ;
        RECT 115.465 102.470 115.625 102.580 ;
        RECT 119.145 102.425 119.315 102.615 ;
        RECT 119.605 102.425 119.775 102.615 ;
        RECT 124.665 102.445 124.835 102.635 ;
        RECT 126.035 102.615 126.205 102.635 ;
        RECT 126.035 102.445 126.215 102.615 ;
        RECT 126.045 102.425 126.215 102.445 ;
        RECT 127.425 102.425 127.595 102.635 ;
        RECT 14.585 101.615 15.955 102.425 ;
        RECT 15.965 101.615 18.715 102.425 ;
        RECT 18.725 101.615 24.235 102.425 ;
        RECT 24.255 101.555 24.685 102.340 ;
        RECT 24.905 101.745 35.275 102.425 ;
        RECT 24.905 101.515 27.115 101.745 ;
        RECT 29.835 101.525 30.765 101.745 ;
        RECT 35.285 101.615 37.115 102.425 ;
        RECT 37.135 101.555 37.565 102.340 ;
        RECT 37.585 101.615 38.955 102.425 ;
        RECT 38.965 101.615 44.475 102.425 ;
        RECT 44.485 101.615 49.995 102.425 ;
        RECT 50.015 101.555 50.445 102.340 ;
        RECT 50.465 101.615 51.835 102.425 ;
        RECT 51.845 101.615 57.355 102.425 ;
        RECT 57.365 101.615 62.875 102.425 ;
        RECT 62.895 101.555 63.325 102.340 ;
        RECT 63.345 101.615 64.715 102.425 ;
        RECT 64.725 101.615 70.235 102.425 ;
        RECT 70.245 101.615 75.755 102.425 ;
        RECT 75.775 101.555 76.205 102.340 ;
        RECT 76.225 101.615 77.595 102.425 ;
        RECT 77.605 101.615 83.115 102.425 ;
        RECT 83.125 101.615 88.635 102.425 ;
        RECT 88.655 101.555 89.085 102.340 ;
        RECT 89.105 101.615 90.935 102.425 ;
        RECT 91.145 101.745 101.515 102.425 ;
        RECT 91.145 101.515 93.355 101.745 ;
        RECT 96.075 101.525 97.005 101.745 ;
        RECT 101.535 101.555 101.965 102.340 ;
        RECT 101.985 101.615 103.355 102.425 ;
        RECT 103.365 101.615 108.875 102.425 ;
        RECT 108.885 101.615 114.395 102.425 ;
        RECT 114.415 101.555 114.845 102.340 ;
        RECT 115.785 101.615 119.455 102.425 ;
        RECT 119.475 101.515 120.825 102.425 ;
        RECT 120.845 101.615 126.355 102.425 ;
        RECT 126.365 101.615 127.735 102.425 ;
      LAYER nwell ;
        RECT 14.390 99.620 127.930 101.225 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.580 211.245 127.740 211.415 ;
        RECT 14.665 210.495 15.875 211.245 ;
        RECT 14.665 209.955 15.185 210.495 ;
        RECT 16.045 210.475 18.635 211.245 ;
        RECT 18.810 210.700 24.155 211.245 ;
        RECT 15.355 209.785 15.875 210.325 ;
        RECT 14.665 208.695 15.875 209.785 ;
        RECT 16.045 209.785 17.255 210.305 ;
        RECT 17.425 209.955 18.635 210.475 ;
        RECT 16.045 208.695 18.635 209.785 ;
        RECT 20.400 209.130 20.750 210.380 ;
        RECT 22.230 209.870 22.570 210.700 ;
        RECT 24.325 210.520 24.615 211.245 ;
        RECT 24.785 210.495 25.995 211.245 ;
        RECT 26.170 210.700 31.515 211.245 ;
        RECT 31.690 210.700 37.035 211.245 ;
        RECT 18.810 208.695 24.155 209.130 ;
        RECT 24.325 208.695 24.615 209.860 ;
        RECT 24.785 209.785 25.305 210.325 ;
        RECT 25.475 209.955 25.995 210.495 ;
        RECT 24.785 208.695 25.995 209.785 ;
        RECT 27.760 209.130 28.110 210.380 ;
        RECT 29.590 209.870 29.930 210.700 ;
        RECT 33.280 209.130 33.630 210.380 ;
        RECT 35.110 209.870 35.450 210.700 ;
        RECT 37.205 210.520 37.495 211.245 ;
        RECT 37.665 210.495 38.875 211.245 ;
        RECT 39.050 210.700 44.395 211.245 ;
        RECT 44.570 210.700 49.915 211.245 ;
        RECT 26.170 208.695 31.515 209.130 ;
        RECT 31.690 208.695 37.035 209.130 ;
        RECT 37.205 208.695 37.495 209.860 ;
        RECT 37.665 209.785 38.185 210.325 ;
        RECT 38.355 209.955 38.875 210.495 ;
        RECT 37.665 208.695 38.875 209.785 ;
        RECT 40.640 209.130 40.990 210.380 ;
        RECT 42.470 209.870 42.810 210.700 ;
        RECT 46.160 209.130 46.510 210.380 ;
        RECT 47.990 209.870 48.330 210.700 ;
        RECT 50.085 210.520 50.375 211.245 ;
        RECT 50.545 210.495 51.755 211.245 ;
        RECT 51.930 210.700 57.275 211.245 ;
        RECT 57.450 210.700 62.795 211.245 ;
        RECT 39.050 208.695 44.395 209.130 ;
        RECT 44.570 208.695 49.915 209.130 ;
        RECT 50.085 208.695 50.375 209.860 ;
        RECT 50.545 209.785 51.065 210.325 ;
        RECT 51.235 209.955 51.755 210.495 ;
        RECT 50.545 208.695 51.755 209.785 ;
        RECT 53.520 209.130 53.870 210.380 ;
        RECT 55.350 209.870 55.690 210.700 ;
        RECT 59.040 209.130 59.390 210.380 ;
        RECT 60.870 209.870 61.210 210.700 ;
        RECT 62.965 210.520 63.255 211.245 ;
        RECT 63.425 210.495 64.635 211.245 ;
        RECT 64.810 210.700 70.155 211.245 ;
        RECT 70.330 210.700 75.675 211.245 ;
        RECT 51.930 208.695 57.275 209.130 ;
        RECT 57.450 208.695 62.795 209.130 ;
        RECT 62.965 208.695 63.255 209.860 ;
        RECT 63.425 209.785 63.945 210.325 ;
        RECT 64.115 209.955 64.635 210.495 ;
        RECT 63.425 208.695 64.635 209.785 ;
        RECT 66.400 209.130 66.750 210.380 ;
        RECT 68.230 209.870 68.570 210.700 ;
        RECT 71.920 209.130 72.270 210.380 ;
        RECT 73.750 209.870 74.090 210.700 ;
        RECT 75.845 210.520 76.135 211.245 ;
        RECT 76.305 210.495 77.515 211.245 ;
        RECT 77.690 210.700 83.035 211.245 ;
        RECT 83.210 210.700 88.555 211.245 ;
        RECT 64.810 208.695 70.155 209.130 ;
        RECT 70.330 208.695 75.675 209.130 ;
        RECT 75.845 208.695 76.135 209.860 ;
        RECT 76.305 209.785 76.825 210.325 ;
        RECT 76.995 209.955 77.515 210.495 ;
        RECT 76.305 208.695 77.515 209.785 ;
        RECT 79.280 209.130 79.630 210.380 ;
        RECT 81.110 209.870 81.450 210.700 ;
        RECT 84.800 209.130 85.150 210.380 ;
        RECT 86.630 209.870 86.970 210.700 ;
        RECT 88.725 210.520 89.015 211.245 ;
        RECT 89.185 210.495 90.395 211.245 ;
        RECT 90.570 210.700 95.915 211.245 ;
        RECT 96.090 210.700 101.435 211.245 ;
        RECT 77.690 208.695 83.035 209.130 ;
        RECT 83.210 208.695 88.555 209.130 ;
        RECT 88.725 208.695 89.015 209.860 ;
        RECT 89.185 209.785 89.705 210.325 ;
        RECT 89.875 209.955 90.395 210.495 ;
        RECT 89.185 208.695 90.395 209.785 ;
        RECT 92.160 209.130 92.510 210.380 ;
        RECT 93.990 209.870 94.330 210.700 ;
        RECT 97.680 209.130 98.030 210.380 ;
        RECT 99.510 209.870 99.850 210.700 ;
        RECT 101.605 210.520 101.895 211.245 ;
        RECT 102.065 210.495 103.275 211.245 ;
        RECT 103.450 210.700 108.795 211.245 ;
        RECT 108.970 210.700 114.315 211.245 ;
        RECT 90.570 208.695 95.915 209.130 ;
        RECT 96.090 208.695 101.435 209.130 ;
        RECT 101.605 208.695 101.895 209.860 ;
        RECT 102.065 209.785 102.585 210.325 ;
        RECT 102.755 209.955 103.275 210.495 ;
        RECT 102.065 208.695 103.275 209.785 ;
        RECT 105.040 209.130 105.390 210.380 ;
        RECT 106.870 209.870 107.210 210.700 ;
        RECT 110.560 209.130 110.910 210.380 ;
        RECT 112.390 209.870 112.730 210.700 ;
        RECT 114.485 210.520 114.775 211.245 ;
        RECT 115.410 210.700 120.755 211.245 ;
        RECT 120.930 210.700 126.275 211.245 ;
        RECT 103.450 208.695 108.795 209.130 ;
        RECT 108.970 208.695 114.315 209.130 ;
        RECT 114.485 208.695 114.775 209.860 ;
        RECT 117.000 209.130 117.350 210.380 ;
        RECT 118.830 209.870 119.170 210.700 ;
        RECT 122.520 209.130 122.870 210.380 ;
        RECT 124.350 209.870 124.690 210.700 ;
        RECT 126.445 210.495 127.655 211.245 ;
        RECT 126.445 209.785 126.965 210.325 ;
        RECT 127.135 209.955 127.655 210.495 ;
        RECT 115.410 208.695 120.755 209.130 ;
        RECT 120.930 208.695 126.275 209.130 ;
        RECT 126.445 208.695 127.655 209.785 ;
        RECT 14.580 208.525 127.740 208.695 ;
        RECT 14.665 207.435 15.875 208.525 ;
        RECT 14.665 206.725 15.185 207.265 ;
        RECT 15.355 206.895 15.875 207.435 ;
        RECT 16.045 207.435 18.635 208.525 ;
        RECT 18.810 208.090 24.155 208.525 ;
        RECT 16.045 206.915 17.255 207.435 ;
        RECT 17.425 206.745 18.635 207.265 ;
        RECT 20.400 206.840 20.750 208.090 ;
        RECT 24.325 207.360 24.615 208.525 ;
        RECT 25.245 207.435 27.835 208.525 ;
        RECT 28.010 208.090 33.355 208.525 ;
        RECT 33.530 208.090 38.875 208.525 ;
        RECT 39.050 208.090 44.395 208.525 ;
        RECT 44.570 208.090 49.915 208.525 ;
        RECT 14.665 205.975 15.875 206.725 ;
        RECT 16.045 205.975 18.635 206.745 ;
        RECT 22.230 206.520 22.570 207.350 ;
        RECT 25.245 206.915 26.455 207.435 ;
        RECT 26.625 206.745 27.835 207.265 ;
        RECT 29.600 206.840 29.950 208.090 ;
        RECT 18.810 205.975 24.155 206.520 ;
        RECT 24.325 205.975 24.615 206.700 ;
        RECT 25.245 205.975 27.835 206.745 ;
        RECT 31.430 206.520 31.770 207.350 ;
        RECT 35.120 206.840 35.470 208.090 ;
        RECT 36.950 206.520 37.290 207.350 ;
        RECT 40.640 206.840 40.990 208.090 ;
        RECT 42.470 206.520 42.810 207.350 ;
        RECT 46.160 206.840 46.510 208.090 ;
        RECT 50.085 207.360 50.375 208.525 ;
        RECT 50.550 208.090 55.895 208.525 ;
        RECT 56.070 208.090 61.415 208.525 ;
        RECT 61.590 208.090 66.935 208.525 ;
        RECT 67.110 208.090 72.455 208.525 ;
        RECT 47.990 206.520 48.330 207.350 ;
        RECT 52.140 206.840 52.490 208.090 ;
        RECT 28.010 205.975 33.355 206.520 ;
        RECT 33.530 205.975 38.875 206.520 ;
        RECT 39.050 205.975 44.395 206.520 ;
        RECT 44.570 205.975 49.915 206.520 ;
        RECT 50.085 205.975 50.375 206.700 ;
        RECT 53.970 206.520 54.310 207.350 ;
        RECT 57.660 206.840 58.010 208.090 ;
        RECT 59.490 206.520 59.830 207.350 ;
        RECT 63.180 206.840 63.530 208.090 ;
        RECT 65.010 206.520 65.350 207.350 ;
        RECT 68.700 206.840 69.050 208.090 ;
        RECT 72.665 207.385 72.895 208.525 ;
        RECT 73.065 207.375 73.395 208.355 ;
        RECT 73.565 207.385 73.775 208.525 ;
        RECT 74.095 207.595 74.265 208.355 ;
        RECT 74.480 207.765 74.810 208.525 ;
        RECT 74.095 207.425 74.810 207.595 ;
        RECT 74.980 207.450 75.235 208.355 ;
        RECT 70.530 206.520 70.870 207.350 ;
        RECT 72.645 206.965 72.975 207.215 ;
        RECT 50.550 205.975 55.895 206.520 ;
        RECT 56.070 205.975 61.415 206.520 ;
        RECT 61.590 205.975 66.935 206.520 ;
        RECT 67.110 205.975 72.455 206.520 ;
        RECT 72.665 205.975 72.895 206.795 ;
        RECT 73.145 206.775 73.395 207.375 ;
        RECT 74.005 206.875 74.360 207.245 ;
        RECT 74.640 207.215 74.810 207.425 ;
        RECT 74.640 206.885 74.895 207.215 ;
        RECT 73.065 206.145 73.395 206.775 ;
        RECT 73.565 205.975 73.775 206.795 ;
        RECT 74.640 206.695 74.810 206.885 ;
        RECT 75.065 206.720 75.235 207.450 ;
        RECT 75.410 207.375 75.670 208.525 ;
        RECT 75.845 207.360 76.135 208.525 ;
        RECT 77.245 208.015 77.545 208.525 ;
        RECT 77.715 208.015 78.095 208.185 ;
        RECT 78.675 208.015 79.305 208.525 ;
        RECT 77.715 207.845 77.885 208.015 ;
        RECT 79.475 207.845 79.805 208.355 ;
        RECT 79.975 208.015 80.275 208.525 ;
        RECT 77.225 207.645 77.885 207.845 ;
        RECT 78.055 207.675 80.275 207.845 ;
        RECT 74.095 206.525 74.810 206.695 ;
        RECT 74.095 206.145 74.265 206.525 ;
        RECT 74.480 205.975 74.810 206.355 ;
        RECT 74.980 206.145 75.235 206.720 ;
        RECT 75.410 205.975 75.670 206.815 ;
        RECT 77.225 206.715 77.395 207.645 ;
        RECT 78.055 207.475 78.225 207.675 ;
        RECT 77.565 207.305 78.225 207.475 ;
        RECT 78.395 207.335 79.935 207.505 ;
        RECT 77.565 206.885 77.735 207.305 ;
        RECT 78.395 207.135 78.565 207.335 ;
        RECT 77.965 206.965 78.565 207.135 ;
        RECT 78.735 206.965 79.430 207.165 ;
        RECT 79.690 206.885 79.935 207.335 ;
        RECT 78.055 206.715 78.965 206.795 ;
        RECT 75.845 205.975 76.135 206.700 ;
        RECT 77.225 206.235 77.545 206.715 ;
        RECT 77.715 206.625 78.965 206.715 ;
        RECT 77.715 206.545 78.225 206.625 ;
        RECT 77.715 206.145 77.945 206.545 ;
        RECT 78.115 205.975 78.465 206.365 ;
        RECT 78.635 206.145 78.965 206.625 ;
        RECT 79.135 205.975 79.305 206.795 ;
        RECT 80.105 206.715 80.275 207.675 ;
        RECT 81.365 207.435 84.875 208.525 ;
        RECT 85.050 208.090 90.395 208.525 ;
        RECT 90.570 208.090 95.915 208.525 ;
        RECT 96.090 208.090 101.435 208.525 ;
        RECT 81.365 206.915 83.055 207.435 ;
        RECT 83.225 206.745 84.875 207.265 ;
        RECT 86.640 206.840 86.990 208.090 ;
        RECT 79.810 206.170 80.275 206.715 ;
        RECT 81.365 205.975 84.875 206.745 ;
        RECT 88.470 206.520 88.810 207.350 ;
        RECT 92.160 206.840 92.510 208.090 ;
        RECT 93.990 206.520 94.330 207.350 ;
        RECT 97.680 206.840 98.030 208.090 ;
        RECT 101.605 207.360 101.895 208.525 ;
        RECT 102.525 207.435 104.195 208.525 ;
        RECT 104.370 208.090 109.715 208.525 ;
        RECT 109.890 208.090 115.235 208.525 ;
        RECT 115.410 208.090 120.755 208.525 ;
        RECT 120.930 208.090 126.275 208.525 ;
        RECT 99.510 206.520 99.850 207.350 ;
        RECT 102.525 206.915 103.275 207.435 ;
        RECT 103.445 206.745 104.195 207.265 ;
        RECT 105.960 206.840 106.310 208.090 ;
        RECT 85.050 205.975 90.395 206.520 ;
        RECT 90.570 205.975 95.915 206.520 ;
        RECT 96.090 205.975 101.435 206.520 ;
        RECT 101.605 205.975 101.895 206.700 ;
        RECT 102.525 205.975 104.195 206.745 ;
        RECT 107.790 206.520 108.130 207.350 ;
        RECT 111.480 206.840 111.830 208.090 ;
        RECT 113.310 206.520 113.650 207.350 ;
        RECT 117.000 206.840 117.350 208.090 ;
        RECT 118.830 206.520 119.170 207.350 ;
        RECT 122.520 206.840 122.870 208.090 ;
        RECT 126.445 207.435 127.655 208.525 ;
        RECT 124.350 206.520 124.690 207.350 ;
        RECT 126.445 206.895 126.965 207.435 ;
        RECT 127.135 206.725 127.655 207.265 ;
        RECT 104.370 205.975 109.715 206.520 ;
        RECT 109.890 205.975 115.235 206.520 ;
        RECT 115.410 205.975 120.755 206.520 ;
        RECT 120.930 205.975 126.275 206.520 ;
        RECT 126.445 205.975 127.655 206.725 ;
        RECT 14.580 205.805 127.740 205.975 ;
        RECT 14.665 205.055 15.875 205.805 ;
        RECT 14.665 204.515 15.185 205.055 ;
        RECT 16.965 205.035 20.475 205.805 ;
        RECT 20.650 205.260 25.995 205.805 ;
        RECT 26.170 205.260 31.515 205.805 ;
        RECT 31.690 205.260 37.035 205.805 ;
        RECT 15.355 204.345 15.875 204.885 ;
        RECT 14.665 203.255 15.875 204.345 ;
        RECT 16.965 204.345 18.655 204.865 ;
        RECT 18.825 204.515 20.475 205.035 ;
        RECT 16.965 203.255 20.475 204.345 ;
        RECT 22.240 203.690 22.590 204.940 ;
        RECT 24.070 204.430 24.410 205.260 ;
        RECT 27.760 203.690 28.110 204.940 ;
        RECT 29.590 204.430 29.930 205.260 ;
        RECT 33.280 203.690 33.630 204.940 ;
        RECT 35.110 204.430 35.450 205.260 ;
        RECT 37.205 205.080 37.495 205.805 ;
        RECT 38.125 205.035 40.715 205.805 ;
        RECT 40.890 205.260 46.235 205.805 ;
        RECT 46.410 205.260 51.755 205.805 ;
        RECT 51.930 205.260 57.275 205.805 ;
        RECT 57.450 205.260 62.795 205.805 ;
        RECT 20.650 203.255 25.995 203.690 ;
        RECT 26.170 203.255 31.515 203.690 ;
        RECT 31.690 203.255 37.035 203.690 ;
        RECT 37.205 203.255 37.495 204.420 ;
        RECT 38.125 204.345 39.335 204.865 ;
        RECT 39.505 204.515 40.715 205.035 ;
        RECT 38.125 203.255 40.715 204.345 ;
        RECT 42.480 203.690 42.830 204.940 ;
        RECT 44.310 204.430 44.650 205.260 ;
        RECT 48.000 203.690 48.350 204.940 ;
        RECT 49.830 204.430 50.170 205.260 ;
        RECT 53.520 203.690 53.870 204.940 ;
        RECT 55.350 204.430 55.690 205.260 ;
        RECT 59.040 203.690 59.390 204.940 ;
        RECT 60.870 204.430 61.210 205.260 ;
        RECT 62.965 205.080 63.255 205.805 ;
        RECT 63.425 205.055 64.635 205.805 ;
        RECT 40.890 203.255 46.235 203.690 ;
        RECT 46.410 203.255 51.755 203.690 ;
        RECT 51.930 203.255 57.275 203.690 ;
        RECT 57.450 203.255 62.795 203.690 ;
        RECT 62.965 203.255 63.255 204.420 ;
        RECT 63.425 204.345 63.945 204.885 ;
        RECT 64.115 204.515 64.635 205.055 ;
        RECT 64.865 204.985 65.075 205.805 ;
        RECT 65.245 205.005 65.575 205.635 ;
        RECT 65.245 204.405 65.495 205.005 ;
        RECT 65.745 204.985 65.975 205.805 ;
        RECT 67.145 204.985 67.375 205.805 ;
        RECT 67.545 205.005 67.875 205.635 ;
        RECT 65.665 204.565 65.995 204.815 ;
        RECT 67.125 204.565 67.455 204.815 ;
        RECT 67.625 204.405 67.875 205.005 ;
        RECT 68.045 204.985 68.255 205.805 ;
        RECT 68.490 205.095 68.745 205.625 ;
        RECT 68.915 205.345 69.220 205.805 ;
        RECT 69.465 205.425 70.535 205.595 ;
        RECT 63.425 203.255 64.635 204.345 ;
        RECT 64.865 203.255 65.075 204.395 ;
        RECT 65.245 203.425 65.575 204.405 ;
        RECT 65.745 203.255 65.975 204.395 ;
        RECT 67.145 203.255 67.375 204.395 ;
        RECT 67.545 203.425 67.875 204.405 ;
        RECT 68.490 204.445 68.700 205.095 ;
        RECT 69.465 205.070 69.785 205.425 ;
        RECT 69.460 204.895 69.785 205.070 ;
        RECT 68.870 204.595 69.785 204.895 ;
        RECT 69.955 204.855 70.195 205.255 ;
        RECT 70.365 205.195 70.535 205.425 ;
        RECT 70.705 205.365 70.895 205.805 ;
        RECT 71.065 205.355 72.015 205.635 ;
        RECT 72.235 205.445 72.585 205.615 ;
        RECT 70.365 205.025 70.895 205.195 ;
        RECT 68.870 204.565 69.610 204.595 ;
        RECT 68.045 203.255 68.255 204.395 ;
        RECT 68.490 203.565 68.745 204.445 ;
        RECT 68.915 203.255 69.220 204.395 ;
        RECT 69.440 203.975 69.610 204.565 ;
        RECT 69.955 204.485 70.495 204.855 ;
        RECT 70.675 204.745 70.895 205.025 ;
        RECT 71.065 204.575 71.235 205.355 ;
        RECT 70.830 204.405 71.235 204.575 ;
        RECT 71.405 204.565 71.755 205.185 ;
        RECT 70.830 204.315 71.000 204.405 ;
        RECT 71.925 204.395 72.135 205.185 ;
        RECT 69.780 204.145 71.000 204.315 ;
        RECT 71.460 204.235 72.135 204.395 ;
        RECT 69.440 203.805 70.240 203.975 ;
        RECT 69.560 203.255 69.890 203.635 ;
        RECT 70.070 203.515 70.240 203.805 ;
        RECT 70.830 203.765 71.000 204.145 ;
        RECT 71.170 204.225 72.135 204.235 ;
        RECT 72.325 205.055 72.585 205.445 ;
        RECT 72.795 205.345 73.125 205.805 ;
        RECT 74.000 205.415 74.855 205.585 ;
        RECT 75.060 205.415 75.555 205.585 ;
        RECT 75.725 205.445 76.055 205.805 ;
        RECT 72.325 204.365 72.495 205.055 ;
        RECT 72.665 204.705 72.835 204.885 ;
        RECT 73.005 204.875 73.795 205.125 ;
        RECT 74.000 204.705 74.170 205.415 ;
        RECT 74.340 204.905 74.695 205.125 ;
        RECT 72.665 204.535 74.355 204.705 ;
        RECT 71.170 203.935 71.630 204.225 ;
        RECT 72.325 204.195 73.825 204.365 ;
        RECT 72.325 204.055 72.495 204.195 ;
        RECT 71.935 203.885 72.495 204.055 ;
        RECT 70.410 203.255 70.660 203.715 ;
        RECT 70.830 203.425 71.700 203.765 ;
        RECT 71.935 203.425 72.105 203.885 ;
        RECT 72.940 203.855 74.015 204.025 ;
        RECT 72.275 203.255 72.645 203.715 ;
        RECT 72.940 203.515 73.110 203.855 ;
        RECT 73.280 203.255 73.610 203.685 ;
        RECT 73.845 203.515 74.015 203.855 ;
        RECT 74.185 203.755 74.355 204.535 ;
        RECT 74.525 204.315 74.695 204.905 ;
        RECT 74.865 204.505 75.215 205.125 ;
        RECT 74.525 203.925 74.990 204.315 ;
        RECT 75.385 204.055 75.555 205.415 ;
        RECT 75.725 204.225 76.185 205.275 ;
        RECT 75.160 203.885 75.555 204.055 ;
        RECT 75.160 203.755 75.330 203.885 ;
        RECT 74.185 203.425 74.865 203.755 ;
        RECT 75.080 203.425 75.330 203.755 ;
        RECT 75.500 203.255 75.750 203.715 ;
        RECT 75.920 203.440 76.245 204.225 ;
        RECT 76.415 203.425 76.585 205.545 ;
        RECT 76.755 205.425 77.085 205.805 ;
        RECT 77.255 205.255 77.510 205.545 ;
        RECT 76.760 205.085 77.510 205.255 ;
        RECT 77.690 205.095 77.945 205.625 ;
        RECT 78.115 205.345 78.420 205.805 ;
        RECT 78.665 205.425 79.735 205.595 ;
        RECT 76.760 204.095 76.990 205.085 ;
        RECT 77.160 204.265 77.510 204.915 ;
        RECT 77.690 204.445 77.900 205.095 ;
        RECT 78.665 205.070 78.985 205.425 ;
        RECT 78.660 204.895 78.985 205.070 ;
        RECT 78.070 204.595 78.985 204.895 ;
        RECT 79.155 204.855 79.395 205.255 ;
        RECT 79.565 205.195 79.735 205.425 ;
        RECT 79.905 205.365 80.095 205.805 ;
        RECT 80.265 205.355 81.215 205.635 ;
        RECT 81.435 205.445 81.785 205.615 ;
        RECT 79.565 205.025 80.095 205.195 ;
        RECT 78.070 204.565 78.810 204.595 ;
        RECT 76.760 203.925 77.510 204.095 ;
        RECT 76.755 203.255 77.085 203.755 ;
        RECT 77.255 203.425 77.510 203.925 ;
        RECT 77.690 203.565 77.945 204.445 ;
        RECT 78.115 203.255 78.420 204.395 ;
        RECT 78.640 203.975 78.810 204.565 ;
        RECT 79.155 204.485 79.695 204.855 ;
        RECT 79.875 204.745 80.095 205.025 ;
        RECT 80.265 204.575 80.435 205.355 ;
        RECT 80.030 204.405 80.435 204.575 ;
        RECT 80.605 204.565 80.955 205.185 ;
        RECT 80.030 204.315 80.200 204.405 ;
        RECT 81.125 204.395 81.335 205.185 ;
        RECT 78.980 204.145 80.200 204.315 ;
        RECT 80.660 204.235 81.335 204.395 ;
        RECT 78.640 203.805 79.440 203.975 ;
        RECT 78.760 203.255 79.090 203.635 ;
        RECT 79.270 203.515 79.440 203.805 ;
        RECT 80.030 203.765 80.200 204.145 ;
        RECT 80.370 204.225 81.335 204.235 ;
        RECT 81.525 205.055 81.785 205.445 ;
        RECT 81.995 205.345 82.325 205.805 ;
        RECT 83.200 205.415 84.055 205.585 ;
        RECT 84.260 205.415 84.755 205.585 ;
        RECT 84.925 205.445 85.255 205.805 ;
        RECT 81.525 204.365 81.695 205.055 ;
        RECT 81.865 204.705 82.035 204.885 ;
        RECT 82.205 204.875 82.995 205.125 ;
        RECT 83.200 204.705 83.370 205.415 ;
        RECT 83.540 204.905 83.895 205.125 ;
        RECT 81.865 204.535 83.555 204.705 ;
        RECT 80.370 203.935 80.830 204.225 ;
        RECT 81.525 204.195 83.025 204.365 ;
        RECT 81.525 204.055 81.695 204.195 ;
        RECT 81.135 203.885 81.695 204.055 ;
        RECT 79.610 203.255 79.860 203.715 ;
        RECT 80.030 203.425 80.900 203.765 ;
        RECT 81.135 203.425 81.305 203.885 ;
        RECT 82.140 203.855 83.215 204.025 ;
        RECT 81.475 203.255 81.845 203.715 ;
        RECT 82.140 203.515 82.310 203.855 ;
        RECT 82.480 203.255 82.810 203.685 ;
        RECT 83.045 203.515 83.215 203.855 ;
        RECT 83.385 203.755 83.555 204.535 ;
        RECT 83.725 204.315 83.895 204.905 ;
        RECT 84.065 204.505 84.415 205.125 ;
        RECT 83.725 203.925 84.190 204.315 ;
        RECT 84.585 204.055 84.755 205.415 ;
        RECT 84.925 204.225 85.385 205.275 ;
        RECT 84.360 203.885 84.755 204.055 ;
        RECT 84.360 203.755 84.530 203.885 ;
        RECT 83.385 203.425 84.065 203.755 ;
        RECT 84.280 203.425 84.530 203.755 ;
        RECT 84.700 203.255 84.950 203.715 ;
        RECT 85.120 203.440 85.445 204.225 ;
        RECT 85.615 203.425 85.785 205.545 ;
        RECT 85.955 205.425 86.285 205.805 ;
        RECT 86.455 205.255 86.710 205.545 ;
        RECT 85.960 205.085 86.710 205.255 ;
        RECT 85.960 204.095 86.190 205.085 ;
        RECT 86.885 205.035 88.555 205.805 ;
        RECT 88.725 205.080 89.015 205.805 ;
        RECT 89.645 205.035 92.235 205.805 ;
        RECT 92.410 205.260 97.755 205.805 ;
        RECT 97.930 205.260 103.275 205.805 ;
        RECT 103.450 205.260 108.795 205.805 ;
        RECT 108.970 205.260 114.315 205.805 ;
        RECT 86.360 204.265 86.710 204.915 ;
        RECT 86.885 204.345 87.635 204.865 ;
        RECT 87.805 204.515 88.555 205.035 ;
        RECT 85.960 203.925 86.710 204.095 ;
        RECT 85.955 203.255 86.285 203.755 ;
        RECT 86.455 203.425 86.710 203.925 ;
        RECT 86.885 203.255 88.555 204.345 ;
        RECT 88.725 203.255 89.015 204.420 ;
        RECT 89.645 204.345 90.855 204.865 ;
        RECT 91.025 204.515 92.235 205.035 ;
        RECT 89.645 203.255 92.235 204.345 ;
        RECT 94.000 203.690 94.350 204.940 ;
        RECT 95.830 204.430 96.170 205.260 ;
        RECT 99.520 203.690 99.870 204.940 ;
        RECT 101.350 204.430 101.690 205.260 ;
        RECT 105.040 203.690 105.390 204.940 ;
        RECT 106.870 204.430 107.210 205.260 ;
        RECT 110.560 203.690 110.910 204.940 ;
        RECT 112.390 204.430 112.730 205.260 ;
        RECT 114.485 205.080 114.775 205.805 ;
        RECT 115.410 205.260 120.755 205.805 ;
        RECT 120.930 205.260 126.275 205.805 ;
        RECT 92.410 203.255 97.755 203.690 ;
        RECT 97.930 203.255 103.275 203.690 ;
        RECT 103.450 203.255 108.795 203.690 ;
        RECT 108.970 203.255 114.315 203.690 ;
        RECT 114.485 203.255 114.775 204.420 ;
        RECT 117.000 203.690 117.350 204.940 ;
        RECT 118.830 204.430 119.170 205.260 ;
        RECT 122.520 203.690 122.870 204.940 ;
        RECT 124.350 204.430 124.690 205.260 ;
        RECT 126.445 205.055 127.655 205.805 ;
        RECT 126.445 204.345 126.965 204.885 ;
        RECT 127.135 204.515 127.655 205.055 ;
        RECT 115.410 203.255 120.755 203.690 ;
        RECT 120.930 203.255 126.275 203.690 ;
        RECT 126.445 203.255 127.655 204.345 ;
        RECT 14.580 203.085 127.740 203.255 ;
        RECT 14.665 201.995 15.875 203.085 ;
        RECT 14.665 201.285 15.185 201.825 ;
        RECT 15.355 201.455 15.875 201.995 ;
        RECT 16.045 201.995 18.635 203.085 ;
        RECT 18.810 202.650 24.155 203.085 ;
        RECT 16.045 201.475 17.255 201.995 ;
        RECT 17.425 201.305 18.635 201.825 ;
        RECT 20.400 201.400 20.750 202.650 ;
        RECT 24.325 201.920 24.615 203.085 ;
        RECT 25.245 201.995 27.835 203.085 ;
        RECT 28.010 202.650 33.355 203.085 ;
        RECT 33.530 202.650 38.875 203.085 ;
        RECT 39.050 202.650 44.395 203.085 ;
        RECT 44.570 202.650 49.915 203.085 ;
        RECT 14.665 200.535 15.875 201.285 ;
        RECT 16.045 200.535 18.635 201.305 ;
        RECT 22.230 201.080 22.570 201.910 ;
        RECT 25.245 201.475 26.455 201.995 ;
        RECT 26.625 201.305 27.835 201.825 ;
        RECT 29.600 201.400 29.950 202.650 ;
        RECT 18.810 200.535 24.155 201.080 ;
        RECT 24.325 200.535 24.615 201.260 ;
        RECT 25.245 200.535 27.835 201.305 ;
        RECT 31.430 201.080 31.770 201.910 ;
        RECT 35.120 201.400 35.470 202.650 ;
        RECT 36.950 201.080 37.290 201.910 ;
        RECT 40.640 201.400 40.990 202.650 ;
        RECT 42.470 201.080 42.810 201.910 ;
        RECT 46.160 201.400 46.510 202.650 ;
        RECT 50.085 201.920 50.375 203.085 ;
        RECT 50.545 201.995 54.055 203.085 ;
        RECT 54.230 202.650 59.575 203.085 ;
        RECT 47.990 201.080 48.330 201.910 ;
        RECT 50.545 201.475 52.235 201.995 ;
        RECT 52.405 201.305 54.055 201.825 ;
        RECT 55.820 201.400 56.170 202.650 ;
        RECT 59.750 202.415 60.005 202.915 ;
        RECT 60.175 202.585 60.505 203.085 ;
        RECT 59.750 202.245 60.500 202.415 ;
        RECT 28.010 200.535 33.355 201.080 ;
        RECT 33.530 200.535 38.875 201.080 ;
        RECT 39.050 200.535 44.395 201.080 ;
        RECT 44.570 200.535 49.915 201.080 ;
        RECT 50.085 200.535 50.375 201.260 ;
        RECT 50.545 200.535 54.055 201.305 ;
        RECT 57.650 201.080 57.990 201.910 ;
        RECT 59.750 201.425 60.100 202.075 ;
        RECT 60.270 201.255 60.500 202.245 ;
        RECT 59.750 201.085 60.500 201.255 ;
        RECT 54.230 200.535 59.575 201.080 ;
        RECT 59.750 200.795 60.005 201.085 ;
        RECT 60.175 200.535 60.505 200.915 ;
        RECT 60.675 200.795 60.845 202.915 ;
        RECT 61.015 202.115 61.340 202.900 ;
        RECT 61.510 202.625 61.760 203.085 ;
        RECT 61.930 202.585 62.180 202.915 ;
        RECT 62.395 202.585 63.075 202.915 ;
        RECT 61.930 202.455 62.100 202.585 ;
        RECT 61.705 202.285 62.100 202.455 ;
        RECT 61.075 201.065 61.535 202.115 ;
        RECT 61.705 200.925 61.875 202.285 ;
        RECT 62.270 202.025 62.735 202.415 ;
        RECT 62.045 201.215 62.395 201.835 ;
        RECT 62.565 201.435 62.735 202.025 ;
        RECT 62.905 201.805 63.075 202.585 ;
        RECT 63.245 202.485 63.415 202.825 ;
        RECT 63.650 202.655 63.980 203.085 ;
        RECT 64.150 202.485 64.320 202.825 ;
        RECT 64.615 202.625 64.985 203.085 ;
        RECT 63.245 202.315 64.320 202.485 ;
        RECT 65.155 202.455 65.325 202.915 ;
        RECT 65.560 202.575 66.430 202.915 ;
        RECT 66.600 202.625 66.850 203.085 ;
        RECT 64.765 202.285 65.325 202.455 ;
        RECT 64.765 202.145 64.935 202.285 ;
        RECT 63.435 201.975 64.935 202.145 ;
        RECT 65.630 202.115 66.090 202.405 ;
        RECT 62.905 201.635 64.595 201.805 ;
        RECT 62.565 201.215 62.920 201.435 ;
        RECT 63.090 200.925 63.260 201.635 ;
        RECT 63.465 201.215 64.255 201.465 ;
        RECT 64.425 201.455 64.595 201.635 ;
        RECT 64.765 201.285 64.935 201.975 ;
        RECT 61.205 200.535 61.535 200.895 ;
        RECT 61.705 200.755 62.200 200.925 ;
        RECT 62.405 200.755 63.260 200.925 ;
        RECT 64.135 200.535 64.465 200.995 ;
        RECT 64.675 200.895 64.935 201.285 ;
        RECT 65.125 202.105 66.090 202.115 ;
        RECT 66.260 202.195 66.430 202.575 ;
        RECT 67.020 202.535 67.190 202.825 ;
        RECT 67.370 202.705 67.700 203.085 ;
        RECT 67.020 202.365 67.820 202.535 ;
        RECT 65.125 201.945 65.800 202.105 ;
        RECT 66.260 202.025 67.480 202.195 ;
        RECT 65.125 201.155 65.335 201.945 ;
        RECT 66.260 201.935 66.430 202.025 ;
        RECT 65.505 201.155 65.855 201.775 ;
        RECT 66.025 201.765 66.430 201.935 ;
        RECT 66.025 200.985 66.195 201.765 ;
        RECT 66.365 201.315 66.585 201.595 ;
        RECT 66.765 201.485 67.305 201.855 ;
        RECT 67.650 201.745 67.820 202.365 ;
        RECT 67.995 202.025 68.165 203.085 ;
        RECT 68.375 202.075 68.665 202.915 ;
        RECT 68.835 202.245 69.005 203.085 ;
        RECT 69.215 202.075 69.465 202.915 ;
        RECT 69.675 202.245 69.845 203.085 ;
        RECT 68.375 201.905 70.100 202.075 ;
        RECT 66.365 201.145 66.895 201.315 ;
        RECT 64.675 200.725 65.025 200.895 ;
        RECT 65.245 200.705 66.195 200.985 ;
        RECT 66.365 200.535 66.555 200.975 ;
        RECT 66.725 200.915 66.895 201.145 ;
        RECT 67.065 201.085 67.305 201.485 ;
        RECT 67.475 201.735 67.820 201.745 ;
        RECT 67.475 201.525 69.505 201.735 ;
        RECT 67.475 201.270 67.800 201.525 ;
        RECT 69.690 201.355 70.100 201.905 ;
        RECT 67.475 200.915 67.795 201.270 ;
        RECT 66.725 200.745 67.795 200.915 ;
        RECT 67.995 200.535 68.165 201.345 ;
        RECT 68.335 201.185 70.100 201.355 ;
        RECT 70.325 201.945 70.585 202.915 ;
        RECT 70.780 202.675 71.110 203.085 ;
        RECT 71.310 202.495 71.480 202.915 ;
        RECT 71.695 202.675 72.365 203.085 ;
        RECT 72.600 202.495 72.770 202.915 ;
        RECT 73.075 202.645 73.405 203.085 ;
        RECT 70.755 202.325 72.770 202.495 ;
        RECT 73.575 202.465 73.750 202.915 ;
        RECT 74.010 202.660 74.345 203.085 ;
        RECT 74.515 202.480 74.700 202.885 ;
        RECT 70.325 201.255 70.495 201.945 ;
        RECT 70.755 201.775 70.925 202.325 ;
        RECT 70.665 201.445 70.925 201.775 ;
        RECT 68.335 200.705 68.665 201.185 ;
        RECT 68.835 200.535 69.005 201.005 ;
        RECT 69.175 200.705 69.505 201.185 ;
        RECT 69.675 200.535 69.845 201.005 ;
        RECT 70.325 200.790 70.665 201.255 ;
        RECT 71.095 201.115 71.435 202.145 ;
        RECT 71.625 201.045 71.895 202.145 ;
        RECT 70.330 200.745 70.665 200.790 ;
        RECT 70.835 200.535 71.165 200.915 ;
        RECT 71.625 200.875 71.935 201.045 ;
        RECT 71.625 200.870 71.895 200.875 ;
        RECT 72.120 200.870 72.400 202.145 ;
        RECT 72.600 201.035 72.770 202.325 ;
        RECT 73.120 202.295 73.750 202.465 ;
        RECT 74.035 202.305 74.700 202.480 ;
        RECT 74.905 202.305 75.235 203.085 ;
        RECT 73.120 201.775 73.290 202.295 ;
        RECT 72.940 201.445 73.290 201.775 ;
        RECT 73.470 201.445 73.835 202.125 ;
        RECT 73.120 201.275 73.290 201.445 ;
        RECT 74.035 201.275 74.375 202.305 ;
        RECT 75.405 202.115 75.675 202.885 ;
        RECT 74.545 201.945 75.675 202.115 ;
        RECT 74.545 201.445 74.795 201.945 ;
        RECT 73.120 201.105 73.750 201.275 ;
        RECT 74.035 201.105 74.720 201.275 ;
        RECT 74.975 201.195 75.335 201.775 ;
        RECT 72.600 200.705 72.830 201.035 ;
        RECT 73.075 200.535 73.405 200.915 ;
        RECT 73.575 200.705 73.750 201.105 ;
        RECT 74.010 200.535 74.345 200.935 ;
        RECT 74.515 200.705 74.720 201.105 ;
        RECT 75.505 201.035 75.675 201.945 ;
        RECT 75.845 201.920 76.135 203.085 ;
        RECT 76.765 202.215 77.040 202.915 ;
        RECT 77.210 202.540 77.465 203.085 ;
        RECT 77.635 202.575 78.115 202.915 ;
        RECT 78.290 202.530 78.895 203.085 ;
        RECT 78.280 202.430 78.895 202.530 ;
        RECT 78.280 202.405 78.465 202.430 ;
        RECT 74.930 200.535 75.205 201.015 ;
        RECT 75.415 200.705 75.675 201.035 ;
        RECT 75.845 200.535 76.135 201.260 ;
        RECT 76.765 201.185 76.935 202.215 ;
        RECT 77.210 202.085 77.965 202.335 ;
        RECT 78.135 202.160 78.465 202.405 ;
        RECT 77.210 202.050 77.980 202.085 ;
        RECT 77.210 202.040 77.995 202.050 ;
        RECT 77.105 202.025 78.000 202.040 ;
        RECT 77.105 202.010 78.020 202.025 ;
        RECT 77.105 202.000 78.040 202.010 ;
        RECT 77.105 201.990 78.065 202.000 ;
        RECT 77.105 201.960 78.135 201.990 ;
        RECT 77.105 201.930 78.155 201.960 ;
        RECT 77.105 201.900 78.175 201.930 ;
        RECT 77.105 201.875 78.205 201.900 ;
        RECT 77.105 201.840 78.240 201.875 ;
        RECT 77.105 201.835 78.270 201.840 ;
        RECT 77.105 201.440 77.335 201.835 ;
        RECT 77.880 201.830 78.270 201.835 ;
        RECT 77.905 201.820 78.270 201.830 ;
        RECT 77.920 201.815 78.270 201.820 ;
        RECT 77.935 201.810 78.270 201.815 ;
        RECT 78.635 201.810 78.895 202.260 ;
        RECT 77.935 201.805 78.895 201.810 ;
        RECT 77.945 201.795 78.895 201.805 ;
        RECT 77.955 201.790 78.895 201.795 ;
        RECT 77.965 201.780 78.895 201.790 ;
        RECT 77.970 201.770 78.895 201.780 ;
        RECT 77.975 201.765 78.895 201.770 ;
        RECT 77.985 201.750 78.895 201.765 ;
        RECT 77.990 201.735 78.895 201.750 ;
        RECT 78.000 201.710 78.895 201.735 ;
        RECT 77.505 201.240 77.835 201.665 ;
        RECT 77.585 201.215 77.835 201.240 ;
        RECT 76.765 200.705 77.025 201.185 ;
        RECT 77.195 200.535 77.445 201.075 ;
        RECT 77.615 200.755 77.835 201.215 ;
        RECT 78.005 201.640 78.895 201.710 ;
        RECT 79.530 201.895 79.785 202.775 ;
        RECT 79.955 201.945 80.260 203.085 ;
        RECT 80.600 202.705 80.930 203.085 ;
        RECT 81.110 202.535 81.280 202.825 ;
        RECT 81.450 202.625 81.700 203.085 ;
        RECT 80.480 202.365 81.280 202.535 ;
        RECT 81.870 202.575 82.740 202.915 ;
        RECT 78.005 200.915 78.175 201.640 ;
        RECT 78.345 201.085 78.895 201.470 ;
        RECT 79.530 201.245 79.740 201.895 ;
        RECT 80.480 201.775 80.650 202.365 ;
        RECT 81.870 202.195 82.040 202.575 ;
        RECT 82.975 202.455 83.145 202.915 ;
        RECT 83.315 202.625 83.685 203.085 ;
        RECT 83.980 202.485 84.150 202.825 ;
        RECT 84.320 202.655 84.650 203.085 ;
        RECT 84.885 202.485 85.055 202.825 ;
        RECT 80.820 202.025 82.040 202.195 ;
        RECT 82.210 202.115 82.670 202.405 ;
        RECT 82.975 202.285 83.535 202.455 ;
        RECT 83.980 202.315 85.055 202.485 ;
        RECT 85.225 202.585 85.905 202.915 ;
        RECT 86.120 202.585 86.370 202.915 ;
        RECT 86.540 202.625 86.790 203.085 ;
        RECT 83.365 202.145 83.535 202.285 ;
        RECT 82.210 202.105 83.175 202.115 ;
        RECT 81.870 201.935 82.040 202.025 ;
        RECT 82.500 201.945 83.175 202.105 ;
        RECT 79.910 201.745 80.650 201.775 ;
        RECT 79.910 201.445 80.825 201.745 ;
        RECT 80.500 201.270 80.825 201.445 ;
        RECT 78.005 200.745 78.895 200.915 ;
        RECT 79.530 200.715 79.785 201.245 ;
        RECT 79.955 200.535 80.260 200.995 ;
        RECT 80.505 200.915 80.825 201.270 ;
        RECT 80.995 201.485 81.535 201.855 ;
        RECT 81.870 201.765 82.275 201.935 ;
        RECT 80.995 201.085 81.235 201.485 ;
        RECT 81.715 201.315 81.935 201.595 ;
        RECT 81.405 201.145 81.935 201.315 ;
        RECT 81.405 200.915 81.575 201.145 ;
        RECT 82.105 200.985 82.275 201.765 ;
        RECT 82.445 201.155 82.795 201.775 ;
        RECT 82.965 201.155 83.175 201.945 ;
        RECT 83.365 201.975 84.865 202.145 ;
        RECT 83.365 201.285 83.535 201.975 ;
        RECT 85.225 201.805 85.395 202.585 ;
        RECT 86.200 202.455 86.370 202.585 ;
        RECT 83.705 201.635 85.395 201.805 ;
        RECT 85.565 202.025 86.030 202.415 ;
        RECT 86.200 202.285 86.595 202.455 ;
        RECT 83.705 201.455 83.875 201.635 ;
        RECT 80.505 200.745 81.575 200.915 ;
        RECT 81.745 200.535 81.935 200.975 ;
        RECT 82.105 200.705 83.055 200.985 ;
        RECT 83.365 200.895 83.625 201.285 ;
        RECT 84.045 201.215 84.835 201.465 ;
        RECT 83.275 200.725 83.625 200.895 ;
        RECT 83.835 200.535 84.165 200.995 ;
        RECT 85.040 200.925 85.210 201.635 ;
        RECT 85.565 201.435 85.735 202.025 ;
        RECT 85.380 201.215 85.735 201.435 ;
        RECT 85.905 201.215 86.255 201.835 ;
        RECT 86.425 200.925 86.595 202.285 ;
        RECT 86.960 202.115 87.285 202.900 ;
        RECT 86.765 201.065 87.225 202.115 ;
        RECT 85.040 200.755 85.895 200.925 ;
        RECT 86.100 200.755 86.595 200.925 ;
        RECT 86.765 200.535 87.095 200.895 ;
        RECT 87.455 200.795 87.625 202.915 ;
        RECT 87.795 202.585 88.125 203.085 ;
        RECT 88.295 202.415 88.550 202.915 ;
        RECT 87.800 202.245 88.550 202.415 ;
        RECT 87.800 201.255 88.030 202.245 ;
        RECT 88.200 201.425 88.550 202.075 ;
        RECT 88.725 201.995 90.395 203.085 ;
        RECT 90.570 202.650 95.915 203.085 ;
        RECT 96.090 202.650 101.435 203.085 ;
        RECT 88.725 201.475 89.475 201.995 ;
        RECT 89.645 201.305 90.395 201.825 ;
        RECT 92.160 201.400 92.510 202.650 ;
        RECT 87.800 201.085 88.550 201.255 ;
        RECT 87.795 200.535 88.125 200.915 ;
        RECT 88.295 200.795 88.550 201.085 ;
        RECT 88.725 200.535 90.395 201.305 ;
        RECT 93.990 201.080 94.330 201.910 ;
        RECT 97.680 201.400 98.030 202.650 ;
        RECT 101.605 201.920 101.895 203.085 ;
        RECT 102.525 201.995 104.195 203.085 ;
        RECT 104.370 202.650 109.715 203.085 ;
        RECT 109.890 202.650 115.235 203.085 ;
        RECT 115.410 202.650 120.755 203.085 ;
        RECT 120.930 202.650 126.275 203.085 ;
        RECT 99.510 201.080 99.850 201.910 ;
        RECT 102.525 201.475 103.275 201.995 ;
        RECT 103.445 201.305 104.195 201.825 ;
        RECT 105.960 201.400 106.310 202.650 ;
        RECT 90.570 200.535 95.915 201.080 ;
        RECT 96.090 200.535 101.435 201.080 ;
        RECT 101.605 200.535 101.895 201.260 ;
        RECT 102.525 200.535 104.195 201.305 ;
        RECT 107.790 201.080 108.130 201.910 ;
        RECT 111.480 201.400 111.830 202.650 ;
        RECT 113.310 201.080 113.650 201.910 ;
        RECT 117.000 201.400 117.350 202.650 ;
        RECT 118.830 201.080 119.170 201.910 ;
        RECT 122.520 201.400 122.870 202.650 ;
        RECT 126.445 201.995 127.655 203.085 ;
        RECT 124.350 201.080 124.690 201.910 ;
        RECT 126.445 201.455 126.965 201.995 ;
        RECT 127.135 201.285 127.655 201.825 ;
        RECT 104.370 200.535 109.715 201.080 ;
        RECT 109.890 200.535 115.235 201.080 ;
        RECT 115.410 200.535 120.755 201.080 ;
        RECT 120.930 200.535 126.275 201.080 ;
        RECT 126.445 200.535 127.655 201.285 ;
        RECT 14.580 200.365 127.740 200.535 ;
        RECT 14.665 199.615 15.875 200.365 ;
        RECT 14.665 199.075 15.185 199.615 ;
        RECT 16.965 199.595 20.475 200.365 ;
        RECT 20.650 199.820 25.995 200.365 ;
        RECT 26.170 199.820 31.515 200.365 ;
        RECT 31.690 199.820 37.035 200.365 ;
        RECT 15.355 198.905 15.875 199.445 ;
        RECT 14.665 197.815 15.875 198.905 ;
        RECT 16.965 198.905 18.655 199.425 ;
        RECT 18.825 199.075 20.475 199.595 ;
        RECT 16.965 197.815 20.475 198.905 ;
        RECT 22.240 198.250 22.590 199.500 ;
        RECT 24.070 198.990 24.410 199.820 ;
        RECT 27.760 198.250 28.110 199.500 ;
        RECT 29.590 198.990 29.930 199.820 ;
        RECT 33.280 198.250 33.630 199.500 ;
        RECT 35.110 198.990 35.450 199.820 ;
        RECT 37.205 199.640 37.495 200.365 ;
        RECT 38.125 199.595 40.715 200.365 ;
        RECT 40.890 199.820 46.235 200.365 ;
        RECT 46.410 199.820 51.755 200.365 ;
        RECT 51.930 199.820 57.275 200.365 ;
        RECT 57.450 199.820 62.795 200.365 ;
        RECT 20.650 197.815 25.995 198.250 ;
        RECT 26.170 197.815 31.515 198.250 ;
        RECT 31.690 197.815 37.035 198.250 ;
        RECT 37.205 197.815 37.495 198.980 ;
        RECT 38.125 198.905 39.335 199.425 ;
        RECT 39.505 199.075 40.715 199.595 ;
        RECT 38.125 197.815 40.715 198.905 ;
        RECT 42.480 198.250 42.830 199.500 ;
        RECT 44.310 198.990 44.650 199.820 ;
        RECT 48.000 198.250 48.350 199.500 ;
        RECT 49.830 198.990 50.170 199.820 ;
        RECT 53.520 198.250 53.870 199.500 ;
        RECT 55.350 198.990 55.690 199.820 ;
        RECT 59.040 198.250 59.390 199.500 ;
        RECT 60.870 198.990 61.210 199.820 ;
        RECT 62.965 199.640 63.255 200.365 ;
        RECT 63.885 199.595 67.395 200.365 ;
        RECT 40.890 197.815 46.235 198.250 ;
        RECT 46.410 197.815 51.755 198.250 ;
        RECT 51.930 197.815 57.275 198.250 ;
        RECT 57.450 197.815 62.795 198.250 ;
        RECT 62.965 197.815 63.255 198.980 ;
        RECT 63.885 198.905 65.575 199.425 ;
        RECT 65.745 199.075 67.395 199.595 ;
        RECT 67.565 199.690 67.825 200.195 ;
        RECT 68.005 199.985 68.335 200.365 ;
        RECT 68.515 199.815 68.685 200.195 ;
        RECT 68.950 199.965 69.285 200.365 ;
        RECT 63.885 197.815 67.395 198.905 ;
        RECT 67.565 198.890 67.735 199.690 ;
        RECT 68.020 199.645 68.685 199.815 ;
        RECT 69.455 199.795 69.660 200.195 ;
        RECT 69.870 199.885 70.145 200.365 ;
        RECT 70.355 199.865 70.615 200.195 ;
        RECT 68.020 199.390 68.190 199.645 ;
        RECT 68.975 199.625 69.660 199.795 ;
        RECT 67.905 199.060 68.190 199.390 ;
        RECT 68.425 199.095 68.755 199.465 ;
        RECT 68.020 198.915 68.190 199.060 ;
        RECT 67.565 197.985 67.835 198.890 ;
        RECT 68.020 198.745 68.685 198.915 ;
        RECT 68.005 197.815 68.335 198.575 ;
        RECT 68.515 197.985 68.685 198.745 ;
        RECT 68.975 198.595 69.315 199.625 ;
        RECT 69.485 198.955 69.735 199.455 ;
        RECT 69.915 199.125 70.275 199.705 ;
        RECT 70.445 198.955 70.615 199.865 ;
        RECT 69.485 198.785 70.615 198.955 ;
        RECT 68.975 198.420 69.640 198.595 ;
        RECT 68.950 197.815 69.285 198.240 ;
        RECT 69.455 198.015 69.640 198.420 ;
        RECT 69.845 197.815 70.175 198.595 ;
        RECT 70.345 198.015 70.615 198.785 ;
        RECT 70.785 197.985 71.045 200.195 ;
        RECT 71.215 199.985 71.545 200.365 ;
        RECT 71.755 199.455 71.950 200.030 ;
        RECT 72.220 199.455 72.405 200.035 ;
        RECT 71.215 198.535 71.385 199.455 ;
        RECT 71.695 199.125 71.950 199.455 ;
        RECT 72.175 199.125 72.405 199.455 ;
        RECT 72.655 200.025 74.135 200.195 ;
        RECT 72.655 199.125 72.825 200.025 ;
        RECT 72.995 199.525 73.545 199.855 ;
        RECT 73.735 199.695 74.135 200.025 ;
        RECT 74.315 199.985 74.645 200.365 ;
        RECT 74.955 199.865 75.215 200.195 ;
        RECT 71.755 198.815 71.950 199.125 ;
        RECT 72.220 198.815 72.405 199.125 ;
        RECT 72.995 198.535 73.165 199.525 ;
        RECT 73.735 199.215 73.905 199.695 ;
        RECT 74.485 199.505 74.695 199.685 ;
        RECT 74.075 199.335 74.695 199.505 ;
        RECT 71.215 198.365 73.165 198.535 ;
        RECT 73.335 199.045 73.905 199.215 ;
        RECT 75.045 199.165 75.215 199.865 ;
        RECT 73.335 198.535 73.505 199.045 ;
        RECT 74.085 198.995 75.215 199.165 ;
        RECT 74.085 198.875 74.255 198.995 ;
        RECT 73.675 198.705 74.255 198.875 ;
        RECT 73.335 198.365 74.075 198.535 ;
        RECT 74.525 198.495 74.875 198.825 ;
        RECT 71.215 197.815 71.545 198.195 ;
        RECT 71.970 197.985 72.140 198.365 ;
        RECT 72.400 197.815 72.730 198.195 ;
        RECT 72.925 197.985 73.095 198.365 ;
        RECT 73.305 197.815 73.635 198.195 ;
        RECT 73.885 197.985 74.075 198.365 ;
        RECT 75.045 198.315 75.215 198.995 ;
        RECT 74.315 197.815 74.645 198.195 ;
        RECT 74.955 197.985 75.215 198.315 ;
        RECT 75.385 199.625 75.770 200.195 ;
        RECT 75.940 199.905 76.265 200.365 ;
        RECT 76.785 199.735 77.065 200.195 ;
        RECT 75.385 198.955 75.665 199.625 ;
        RECT 75.940 199.565 77.065 199.735 ;
        RECT 75.940 199.455 76.390 199.565 ;
        RECT 75.835 199.125 76.390 199.455 ;
        RECT 77.255 199.395 77.655 200.195 ;
        RECT 78.055 199.905 78.325 200.365 ;
        RECT 78.495 199.735 78.780 200.195 ;
        RECT 75.385 197.985 75.770 198.955 ;
        RECT 75.940 198.665 76.390 199.125 ;
        RECT 76.560 198.835 77.655 199.395 ;
        RECT 75.940 198.445 77.065 198.665 ;
        RECT 75.940 197.815 76.265 198.275 ;
        RECT 76.785 197.985 77.065 198.445 ;
        RECT 77.255 197.985 77.655 198.835 ;
        RECT 77.825 199.565 78.780 199.735 ;
        RECT 79.100 199.625 79.715 200.195 ;
        RECT 79.885 199.855 80.100 200.365 ;
        RECT 80.330 199.855 80.610 200.185 ;
        RECT 80.790 199.855 81.030 200.365 ;
        RECT 77.825 198.665 78.035 199.565 ;
        RECT 78.205 198.835 78.895 199.395 ;
        RECT 77.825 198.445 78.780 198.665 ;
        RECT 78.055 197.815 78.325 198.275 ;
        RECT 78.495 197.985 78.780 198.445 ;
        RECT 79.100 198.605 79.415 199.625 ;
        RECT 79.585 198.955 79.755 199.455 ;
        RECT 80.005 199.125 80.270 199.685 ;
        RECT 80.440 198.955 80.610 199.855 ;
        RECT 80.780 199.125 81.135 199.685 ;
        RECT 81.365 199.565 82.060 200.195 ;
        RECT 82.265 199.565 82.575 200.365 ;
        RECT 82.835 199.815 83.005 200.195 ;
        RECT 83.185 199.985 83.515 200.365 ;
        RECT 82.835 199.645 83.500 199.815 ;
        RECT 83.695 199.690 83.955 200.195 ;
        RECT 81.385 199.125 81.720 199.375 ;
        RECT 81.890 198.965 82.060 199.565 ;
        RECT 82.230 199.125 82.565 199.395 ;
        RECT 82.765 199.095 83.095 199.465 ;
        RECT 83.330 199.390 83.500 199.645 ;
        RECT 83.330 199.060 83.615 199.390 ;
        RECT 79.585 198.785 81.010 198.955 ;
        RECT 79.100 197.985 79.635 198.605 ;
        RECT 79.805 197.815 80.135 198.615 ;
        RECT 80.620 198.610 81.010 198.785 ;
        RECT 81.365 197.815 81.625 198.955 ;
        RECT 81.795 197.985 82.125 198.965 ;
        RECT 82.295 197.815 82.575 198.955 ;
        RECT 83.330 198.915 83.500 199.060 ;
        RECT 82.835 198.745 83.500 198.915 ;
        RECT 83.785 198.890 83.955 199.690 ;
        RECT 84.165 199.545 84.395 200.365 ;
        RECT 84.565 199.565 84.895 200.195 ;
        RECT 84.145 199.125 84.475 199.375 ;
        RECT 84.645 198.965 84.895 199.565 ;
        RECT 85.065 199.545 85.275 200.365 ;
        RECT 85.565 199.545 85.775 200.365 ;
        RECT 85.945 199.565 86.275 200.195 ;
        RECT 82.835 197.985 83.005 198.745 ;
        RECT 83.185 197.815 83.515 198.575 ;
        RECT 83.685 197.985 83.955 198.890 ;
        RECT 84.165 197.815 84.395 198.955 ;
        RECT 84.565 197.985 84.895 198.965 ;
        RECT 85.945 198.965 86.195 199.565 ;
        RECT 86.445 199.545 86.675 200.365 ;
        RECT 86.885 199.595 88.555 200.365 ;
        RECT 88.725 199.640 89.015 200.365 ;
        RECT 89.645 199.595 91.315 200.365 ;
        RECT 91.490 199.820 96.835 200.365 ;
        RECT 86.365 199.125 86.695 199.375 ;
        RECT 85.065 197.815 85.275 198.955 ;
        RECT 85.565 197.815 85.775 198.955 ;
        RECT 85.945 197.985 86.275 198.965 ;
        RECT 86.445 197.815 86.675 198.955 ;
        RECT 86.885 198.905 87.635 199.425 ;
        RECT 87.805 199.075 88.555 199.595 ;
        RECT 86.885 197.815 88.555 198.905 ;
        RECT 88.725 197.815 89.015 198.980 ;
        RECT 89.645 198.905 90.395 199.425 ;
        RECT 90.565 199.075 91.315 199.595 ;
        RECT 89.645 197.815 91.315 198.905 ;
        RECT 93.080 198.250 93.430 199.500 ;
        RECT 94.910 198.990 95.250 199.820 ;
        RECT 97.010 199.655 97.265 200.185 ;
        RECT 97.435 199.905 97.740 200.365 ;
        RECT 97.985 199.985 99.055 200.155 ;
        RECT 97.010 199.005 97.220 199.655 ;
        RECT 97.985 199.630 98.305 199.985 ;
        RECT 97.980 199.455 98.305 199.630 ;
        RECT 97.390 199.155 98.305 199.455 ;
        RECT 98.475 199.415 98.715 199.815 ;
        RECT 98.885 199.755 99.055 199.985 ;
        RECT 99.225 199.925 99.415 200.365 ;
        RECT 99.585 199.915 100.535 200.195 ;
        RECT 100.755 200.005 101.105 200.175 ;
        RECT 98.885 199.585 99.415 199.755 ;
        RECT 97.390 199.125 98.130 199.155 ;
        RECT 91.490 197.815 96.835 198.250 ;
        RECT 97.010 198.125 97.265 199.005 ;
        RECT 97.435 197.815 97.740 198.955 ;
        RECT 97.960 198.535 98.130 199.125 ;
        RECT 98.475 199.045 99.015 199.415 ;
        RECT 99.195 199.305 99.415 199.585 ;
        RECT 99.585 199.135 99.755 199.915 ;
        RECT 99.350 198.965 99.755 199.135 ;
        RECT 99.925 199.125 100.275 199.745 ;
        RECT 99.350 198.875 99.520 198.965 ;
        RECT 100.445 198.955 100.655 199.745 ;
        RECT 98.300 198.705 99.520 198.875 ;
        RECT 99.980 198.795 100.655 198.955 ;
        RECT 97.960 198.365 98.760 198.535 ;
        RECT 98.080 197.815 98.410 198.195 ;
        RECT 98.590 198.075 98.760 198.365 ;
        RECT 99.350 198.325 99.520 198.705 ;
        RECT 99.690 198.785 100.655 198.795 ;
        RECT 100.845 199.615 101.105 200.005 ;
        RECT 101.315 199.905 101.645 200.365 ;
        RECT 102.520 199.975 103.375 200.145 ;
        RECT 103.580 199.975 104.075 200.145 ;
        RECT 104.245 200.005 104.575 200.365 ;
        RECT 100.845 198.925 101.015 199.615 ;
        RECT 101.185 199.265 101.355 199.445 ;
        RECT 101.525 199.435 102.315 199.685 ;
        RECT 102.520 199.265 102.690 199.975 ;
        RECT 102.860 199.465 103.215 199.685 ;
        RECT 101.185 199.095 102.875 199.265 ;
        RECT 99.690 198.495 100.150 198.785 ;
        RECT 100.845 198.755 102.345 198.925 ;
        RECT 100.845 198.615 101.015 198.755 ;
        RECT 100.455 198.445 101.015 198.615 ;
        RECT 98.930 197.815 99.180 198.275 ;
        RECT 99.350 197.985 100.220 198.325 ;
        RECT 100.455 197.985 100.625 198.445 ;
        RECT 101.460 198.415 102.535 198.585 ;
        RECT 100.795 197.815 101.165 198.275 ;
        RECT 101.460 198.075 101.630 198.415 ;
        RECT 101.800 197.815 102.130 198.245 ;
        RECT 102.365 198.075 102.535 198.415 ;
        RECT 102.705 198.315 102.875 199.095 ;
        RECT 103.045 198.875 103.215 199.465 ;
        RECT 103.385 199.065 103.735 199.685 ;
        RECT 103.045 198.485 103.510 198.875 ;
        RECT 103.905 198.615 104.075 199.975 ;
        RECT 104.245 198.785 104.705 199.835 ;
        RECT 103.680 198.445 104.075 198.615 ;
        RECT 103.680 198.315 103.850 198.445 ;
        RECT 102.705 197.985 103.385 198.315 ;
        RECT 103.600 197.985 103.850 198.315 ;
        RECT 104.020 197.815 104.270 198.275 ;
        RECT 104.440 198.000 104.765 198.785 ;
        RECT 104.935 197.985 105.105 200.105 ;
        RECT 105.275 199.985 105.605 200.365 ;
        RECT 105.775 199.815 106.030 200.105 ;
        RECT 105.280 199.645 106.030 199.815 ;
        RECT 105.280 198.655 105.510 199.645 ;
        RECT 106.205 199.595 108.795 200.365 ;
        RECT 108.970 199.820 114.315 200.365 ;
        RECT 105.680 198.825 106.030 199.475 ;
        RECT 106.205 198.905 107.415 199.425 ;
        RECT 107.585 199.075 108.795 199.595 ;
        RECT 105.280 198.485 106.030 198.655 ;
        RECT 105.275 197.815 105.605 198.315 ;
        RECT 105.775 197.985 106.030 198.485 ;
        RECT 106.205 197.815 108.795 198.905 ;
        RECT 110.560 198.250 110.910 199.500 ;
        RECT 112.390 198.990 112.730 199.820 ;
        RECT 114.485 199.640 114.775 200.365 ;
        RECT 115.410 199.820 120.755 200.365 ;
        RECT 120.930 199.820 126.275 200.365 ;
        RECT 108.970 197.815 114.315 198.250 ;
        RECT 114.485 197.815 114.775 198.980 ;
        RECT 117.000 198.250 117.350 199.500 ;
        RECT 118.830 198.990 119.170 199.820 ;
        RECT 122.520 198.250 122.870 199.500 ;
        RECT 124.350 198.990 124.690 199.820 ;
        RECT 126.445 199.615 127.655 200.365 ;
        RECT 126.445 198.905 126.965 199.445 ;
        RECT 127.135 199.075 127.655 199.615 ;
        RECT 115.410 197.815 120.755 198.250 ;
        RECT 120.930 197.815 126.275 198.250 ;
        RECT 126.445 197.815 127.655 198.905 ;
        RECT 14.580 197.645 127.740 197.815 ;
        RECT 14.665 196.555 15.875 197.645 ;
        RECT 14.665 195.845 15.185 196.385 ;
        RECT 15.355 196.015 15.875 196.555 ;
        RECT 16.045 196.555 18.635 197.645 ;
        RECT 18.810 197.210 24.155 197.645 ;
        RECT 16.045 196.035 17.255 196.555 ;
        RECT 17.425 195.865 18.635 196.385 ;
        RECT 20.400 195.960 20.750 197.210 ;
        RECT 24.325 196.480 24.615 197.645 ;
        RECT 25.245 196.555 27.835 197.645 ;
        RECT 28.010 197.210 33.355 197.645 ;
        RECT 33.530 197.210 38.875 197.645 ;
        RECT 39.050 197.210 44.395 197.645 ;
        RECT 44.570 197.210 49.915 197.645 ;
        RECT 14.665 195.095 15.875 195.845 ;
        RECT 16.045 195.095 18.635 195.865 ;
        RECT 22.230 195.640 22.570 196.470 ;
        RECT 25.245 196.035 26.455 196.555 ;
        RECT 26.625 195.865 27.835 196.385 ;
        RECT 29.600 195.960 29.950 197.210 ;
        RECT 18.810 195.095 24.155 195.640 ;
        RECT 24.325 195.095 24.615 195.820 ;
        RECT 25.245 195.095 27.835 195.865 ;
        RECT 31.430 195.640 31.770 196.470 ;
        RECT 35.120 195.960 35.470 197.210 ;
        RECT 36.950 195.640 37.290 196.470 ;
        RECT 40.640 195.960 40.990 197.210 ;
        RECT 42.470 195.640 42.810 196.470 ;
        RECT 46.160 195.960 46.510 197.210 ;
        RECT 50.085 196.480 50.375 197.645 ;
        RECT 51.005 196.555 52.675 197.645 ;
        RECT 47.990 195.640 48.330 196.470 ;
        RECT 51.005 196.035 51.755 196.555 ;
        RECT 52.905 196.505 53.115 197.645 ;
        RECT 53.285 196.495 53.615 197.475 ;
        RECT 53.785 196.505 54.015 197.645 ;
        RECT 54.340 197.015 54.625 197.475 ;
        RECT 54.795 197.185 55.065 197.645 ;
        RECT 54.340 196.795 55.295 197.015 ;
        RECT 51.925 195.865 52.675 196.385 ;
        RECT 28.010 195.095 33.355 195.640 ;
        RECT 33.530 195.095 38.875 195.640 ;
        RECT 39.050 195.095 44.395 195.640 ;
        RECT 44.570 195.095 49.915 195.640 ;
        RECT 50.085 195.095 50.375 195.820 ;
        RECT 51.005 195.095 52.675 195.865 ;
        RECT 52.905 195.095 53.115 195.915 ;
        RECT 53.285 195.895 53.535 196.495 ;
        RECT 53.705 196.085 54.035 196.335 ;
        RECT 54.225 196.065 54.915 196.625 ;
        RECT 53.285 195.265 53.615 195.895 ;
        RECT 53.785 195.095 54.015 195.915 ;
        RECT 55.085 195.895 55.295 196.795 ;
        RECT 54.340 195.725 55.295 195.895 ;
        RECT 55.465 196.625 55.865 197.475 ;
        RECT 56.055 197.015 56.335 197.475 ;
        RECT 56.855 197.185 57.180 197.645 ;
        RECT 56.055 196.795 57.180 197.015 ;
        RECT 55.465 196.065 56.560 196.625 ;
        RECT 56.730 196.335 57.180 196.795 ;
        RECT 57.350 196.505 57.735 197.475 ;
        RECT 57.910 197.210 63.255 197.645 ;
        RECT 63.430 197.210 68.775 197.645 ;
        RECT 54.340 195.265 54.625 195.725 ;
        RECT 54.795 195.095 55.065 195.555 ;
        RECT 55.465 195.265 55.865 196.065 ;
        RECT 56.730 196.005 57.285 196.335 ;
        RECT 56.730 195.895 57.180 196.005 ;
        RECT 56.055 195.725 57.180 195.895 ;
        RECT 57.455 195.835 57.735 196.505 ;
        RECT 59.500 195.960 59.850 197.210 ;
        RECT 56.055 195.265 56.335 195.725 ;
        RECT 56.855 195.095 57.180 195.555 ;
        RECT 57.350 195.265 57.735 195.835 ;
        RECT 61.330 195.640 61.670 196.470 ;
        RECT 65.020 195.960 65.370 197.210 ;
        RECT 68.945 196.775 69.220 197.475 ;
        RECT 69.390 197.100 69.645 197.645 ;
        RECT 69.815 197.135 70.295 197.475 ;
        RECT 70.470 197.090 71.075 197.645 ;
        RECT 70.460 196.990 71.075 197.090 ;
        RECT 70.460 196.965 70.645 196.990 ;
        RECT 66.850 195.640 67.190 196.470 ;
        RECT 68.945 195.745 69.115 196.775 ;
        RECT 69.390 196.645 70.145 196.895 ;
        RECT 70.315 196.720 70.645 196.965 ;
        RECT 69.390 196.610 70.160 196.645 ;
        RECT 69.390 196.600 70.175 196.610 ;
        RECT 69.285 196.585 70.180 196.600 ;
        RECT 69.285 196.570 70.200 196.585 ;
        RECT 69.285 196.560 70.220 196.570 ;
        RECT 69.285 196.550 70.245 196.560 ;
        RECT 69.285 196.520 70.315 196.550 ;
        RECT 69.285 196.490 70.335 196.520 ;
        RECT 69.285 196.460 70.355 196.490 ;
        RECT 69.285 196.435 70.385 196.460 ;
        RECT 69.285 196.400 70.420 196.435 ;
        RECT 69.285 196.395 70.450 196.400 ;
        RECT 69.285 196.000 69.515 196.395 ;
        RECT 70.060 196.390 70.450 196.395 ;
        RECT 70.085 196.380 70.450 196.390 ;
        RECT 70.100 196.375 70.450 196.380 ;
        RECT 70.115 196.370 70.450 196.375 ;
        RECT 70.815 196.370 71.075 196.820 ;
        RECT 70.115 196.365 71.075 196.370 ;
        RECT 70.125 196.355 71.075 196.365 ;
        RECT 70.135 196.350 71.075 196.355 ;
        RECT 70.145 196.340 71.075 196.350 ;
        RECT 70.150 196.330 71.075 196.340 ;
        RECT 70.155 196.325 71.075 196.330 ;
        RECT 70.165 196.310 71.075 196.325 ;
        RECT 70.170 196.295 71.075 196.310 ;
        RECT 70.180 196.270 71.075 196.295 ;
        RECT 69.685 195.800 70.015 196.225 ;
        RECT 57.910 195.095 63.255 195.640 ;
        RECT 63.430 195.095 68.775 195.640 ;
        RECT 68.945 195.265 69.205 195.745 ;
        RECT 69.375 195.095 69.625 195.635 ;
        RECT 69.795 195.315 70.015 195.800 ;
        RECT 70.185 196.200 71.075 196.270 ;
        RECT 71.255 196.585 71.585 197.435 ;
        RECT 70.185 195.475 70.355 196.200 ;
        RECT 70.525 195.645 71.075 196.030 ;
        RECT 71.255 195.820 71.445 196.585 ;
        RECT 71.755 196.505 72.005 197.645 ;
        RECT 72.195 197.005 72.445 197.425 ;
        RECT 72.675 197.175 73.005 197.645 ;
        RECT 73.235 197.005 73.485 197.425 ;
        RECT 72.195 196.835 73.485 197.005 ;
        RECT 73.665 197.005 73.995 197.435 ;
        RECT 73.665 196.835 74.120 197.005 ;
        RECT 72.185 196.335 72.400 196.665 ;
        RECT 71.615 196.005 71.925 196.335 ;
        RECT 72.095 196.005 72.400 196.335 ;
        RECT 72.575 196.005 72.860 196.665 ;
        RECT 73.055 196.005 73.320 196.665 ;
        RECT 73.535 196.005 73.780 196.665 ;
        RECT 71.755 195.835 71.925 196.005 ;
        RECT 73.950 195.835 74.120 196.835 ;
        RECT 74.465 196.555 75.675 197.645 ;
        RECT 74.465 196.015 74.985 196.555 ;
        RECT 75.845 196.480 76.135 197.645 ;
        RECT 76.305 196.555 79.815 197.645 ;
        RECT 79.990 197.210 85.335 197.645 ;
        RECT 75.155 195.845 75.675 196.385 ;
        RECT 76.305 196.035 77.995 196.555 ;
        RECT 78.165 195.865 79.815 196.385 ;
        RECT 81.580 195.960 81.930 197.210 ;
        RECT 85.880 196.665 86.135 197.335 ;
        RECT 86.315 196.845 86.600 197.645 ;
        RECT 86.780 196.925 87.110 197.435 ;
        RECT 70.185 195.305 71.075 195.475 ;
        RECT 71.255 195.310 71.585 195.820 ;
        RECT 71.755 195.665 74.120 195.835 ;
        RECT 71.755 195.095 72.085 195.495 ;
        RECT 73.135 195.325 73.465 195.665 ;
        RECT 73.635 195.095 73.965 195.495 ;
        RECT 74.465 195.095 75.675 195.845 ;
        RECT 75.845 195.095 76.135 195.820 ;
        RECT 76.305 195.095 79.815 195.865 ;
        RECT 83.410 195.640 83.750 196.470 ;
        RECT 85.880 195.805 86.060 196.665 ;
        RECT 86.780 196.335 87.030 196.925 ;
        RECT 87.380 196.775 87.550 197.385 ;
        RECT 87.720 196.955 88.050 197.645 ;
        RECT 88.280 197.095 88.520 197.385 ;
        RECT 88.720 197.265 89.140 197.645 ;
        RECT 89.320 197.175 89.950 197.425 ;
        RECT 90.420 197.265 90.750 197.645 ;
        RECT 89.320 197.095 89.490 197.175 ;
        RECT 90.920 197.095 91.090 197.385 ;
        RECT 91.270 197.265 91.650 197.645 ;
        RECT 91.890 197.260 92.720 197.430 ;
        RECT 88.280 196.925 89.490 197.095 ;
        RECT 86.230 196.005 87.030 196.335 ;
        RECT 79.990 195.095 85.335 195.640 ;
        RECT 85.880 195.605 86.135 195.805 ;
        RECT 85.795 195.435 86.135 195.605 ;
        RECT 85.880 195.275 86.135 195.435 ;
        RECT 86.315 195.095 86.600 195.555 ;
        RECT 86.780 195.355 87.030 196.005 ;
        RECT 87.230 196.755 87.550 196.775 ;
        RECT 87.230 196.585 89.150 196.755 ;
        RECT 87.230 195.690 87.420 196.585 ;
        RECT 89.320 196.415 89.490 196.925 ;
        RECT 89.660 196.665 90.180 196.975 ;
        RECT 87.590 196.245 89.490 196.415 ;
        RECT 87.590 196.185 87.920 196.245 ;
        RECT 88.070 196.015 88.400 196.075 ;
        RECT 87.740 195.745 88.400 196.015 ;
        RECT 87.230 195.360 87.550 195.690 ;
        RECT 87.730 195.095 88.390 195.575 ;
        RECT 88.590 195.485 88.760 196.245 ;
        RECT 89.660 196.075 89.840 196.485 ;
        RECT 88.930 195.905 89.260 196.025 ;
        RECT 90.010 195.905 90.180 196.665 ;
        RECT 88.930 195.735 90.180 195.905 ;
        RECT 90.350 196.845 91.720 197.095 ;
        RECT 90.350 196.075 90.540 196.845 ;
        RECT 91.470 196.585 91.720 196.845 ;
        RECT 90.710 196.415 90.960 196.575 ;
        RECT 91.890 196.415 92.060 197.260 ;
        RECT 92.955 196.975 93.125 197.475 ;
        RECT 93.295 197.145 93.625 197.645 ;
        RECT 92.230 196.585 92.730 196.965 ;
        RECT 92.955 196.805 93.650 196.975 ;
        RECT 90.710 196.245 92.060 196.415 ;
        RECT 91.640 196.205 92.060 196.245 ;
        RECT 90.350 195.735 90.770 196.075 ;
        RECT 91.060 195.745 91.470 196.075 ;
        RECT 88.590 195.315 89.440 195.485 ;
        RECT 90.000 195.095 90.320 195.555 ;
        RECT 90.520 195.305 90.770 195.735 ;
        RECT 91.060 195.095 91.470 195.535 ;
        RECT 91.640 195.475 91.810 196.205 ;
        RECT 91.980 195.655 92.330 196.025 ;
        RECT 92.510 195.715 92.730 196.585 ;
        RECT 92.900 196.015 93.310 196.635 ;
        RECT 93.480 195.835 93.650 196.805 ;
        RECT 92.955 195.645 93.650 195.835 ;
        RECT 91.640 195.275 92.655 195.475 ;
        RECT 92.955 195.315 93.125 195.645 ;
        RECT 93.295 195.095 93.625 195.475 ;
        RECT 93.840 195.355 94.065 197.475 ;
        RECT 94.235 197.145 94.565 197.645 ;
        RECT 94.735 196.975 94.905 197.475 ;
        RECT 94.240 196.805 94.905 196.975 ;
        RECT 94.240 195.815 94.470 196.805 ;
        RECT 94.640 195.985 94.990 196.635 ;
        RECT 95.165 196.555 97.755 197.645 ;
        RECT 98.040 197.015 98.325 197.475 ;
        RECT 98.495 197.185 98.765 197.645 ;
        RECT 98.040 196.795 98.995 197.015 ;
        RECT 95.165 196.035 96.375 196.555 ;
        RECT 96.545 195.865 97.755 196.385 ;
        RECT 97.925 196.065 98.615 196.625 ;
        RECT 98.785 195.895 98.995 196.795 ;
        RECT 94.240 195.645 94.905 195.815 ;
        RECT 94.235 195.095 94.565 195.475 ;
        RECT 94.735 195.355 94.905 195.645 ;
        RECT 95.165 195.095 97.755 195.865 ;
        RECT 98.040 195.725 98.995 195.895 ;
        RECT 99.165 196.625 99.565 197.475 ;
        RECT 99.755 197.015 100.035 197.475 ;
        RECT 100.555 197.185 100.880 197.645 ;
        RECT 99.755 196.795 100.880 197.015 ;
        RECT 99.165 196.065 100.260 196.625 ;
        RECT 100.430 196.335 100.880 196.795 ;
        RECT 101.050 196.505 101.435 197.475 ;
        RECT 98.040 195.265 98.325 195.725 ;
        RECT 98.495 195.095 98.765 195.555 ;
        RECT 99.165 195.265 99.565 196.065 ;
        RECT 100.430 196.005 100.985 196.335 ;
        RECT 100.430 195.895 100.880 196.005 ;
        RECT 99.755 195.725 100.880 195.895 ;
        RECT 101.155 195.835 101.435 196.505 ;
        RECT 101.605 196.480 101.895 197.645 ;
        RECT 102.065 196.555 104.655 197.645 ;
        RECT 104.830 197.210 110.175 197.645 ;
        RECT 102.065 196.035 103.275 196.555 ;
        RECT 103.445 195.865 104.655 196.385 ;
        RECT 106.420 195.960 106.770 197.210 ;
        RECT 99.755 195.265 100.035 195.725 ;
        RECT 100.555 195.095 100.880 195.555 ;
        RECT 101.050 195.265 101.435 195.835 ;
        RECT 101.605 195.095 101.895 195.820 ;
        RECT 102.065 195.095 104.655 195.865 ;
        RECT 108.250 195.640 108.590 196.470 ;
        RECT 110.350 196.455 110.605 197.335 ;
        RECT 110.775 196.505 111.080 197.645 ;
        RECT 111.420 197.265 111.750 197.645 ;
        RECT 111.930 197.095 112.100 197.385 ;
        RECT 112.270 197.185 112.520 197.645 ;
        RECT 111.300 196.925 112.100 197.095 ;
        RECT 112.690 197.135 113.560 197.475 ;
        RECT 110.350 195.805 110.560 196.455 ;
        RECT 111.300 196.335 111.470 196.925 ;
        RECT 112.690 196.755 112.860 197.135 ;
        RECT 113.795 197.015 113.965 197.475 ;
        RECT 114.135 197.185 114.505 197.645 ;
        RECT 114.800 197.045 114.970 197.385 ;
        RECT 115.140 197.215 115.470 197.645 ;
        RECT 115.705 197.045 115.875 197.385 ;
        RECT 111.640 196.585 112.860 196.755 ;
        RECT 113.030 196.675 113.490 196.965 ;
        RECT 113.795 196.845 114.355 197.015 ;
        RECT 114.800 196.875 115.875 197.045 ;
        RECT 116.045 197.145 116.725 197.475 ;
        RECT 116.940 197.145 117.190 197.475 ;
        RECT 117.360 197.185 117.610 197.645 ;
        RECT 114.185 196.705 114.355 196.845 ;
        RECT 113.030 196.665 113.995 196.675 ;
        RECT 112.690 196.495 112.860 196.585 ;
        RECT 113.320 196.505 113.995 196.665 ;
        RECT 110.730 196.305 111.470 196.335 ;
        RECT 110.730 196.005 111.645 196.305 ;
        RECT 111.320 195.830 111.645 196.005 ;
        RECT 104.830 195.095 110.175 195.640 ;
        RECT 110.350 195.275 110.605 195.805 ;
        RECT 110.775 195.095 111.080 195.555 ;
        RECT 111.325 195.475 111.645 195.830 ;
        RECT 111.815 196.045 112.355 196.415 ;
        RECT 112.690 196.325 113.095 196.495 ;
        RECT 111.815 195.645 112.055 196.045 ;
        RECT 112.535 195.875 112.755 196.155 ;
        RECT 112.225 195.705 112.755 195.875 ;
        RECT 112.225 195.475 112.395 195.705 ;
        RECT 112.925 195.545 113.095 196.325 ;
        RECT 113.265 195.715 113.615 196.335 ;
        RECT 113.785 195.715 113.995 196.505 ;
        RECT 114.185 196.535 115.685 196.705 ;
        RECT 114.185 195.845 114.355 196.535 ;
        RECT 116.045 196.365 116.215 197.145 ;
        RECT 117.020 197.015 117.190 197.145 ;
        RECT 114.525 196.195 116.215 196.365 ;
        RECT 116.385 196.585 116.850 196.975 ;
        RECT 117.020 196.845 117.415 197.015 ;
        RECT 114.525 196.015 114.695 196.195 ;
        RECT 111.325 195.305 112.395 195.475 ;
        RECT 112.565 195.095 112.755 195.535 ;
        RECT 112.925 195.265 113.875 195.545 ;
        RECT 114.185 195.455 114.445 195.845 ;
        RECT 114.865 195.775 115.655 196.025 ;
        RECT 114.095 195.285 114.445 195.455 ;
        RECT 114.655 195.095 114.985 195.555 ;
        RECT 115.860 195.485 116.030 196.195 ;
        RECT 116.385 195.995 116.555 196.585 ;
        RECT 116.200 195.775 116.555 195.995 ;
        RECT 116.725 195.775 117.075 196.395 ;
        RECT 117.245 195.485 117.415 196.845 ;
        RECT 117.780 196.675 118.105 197.460 ;
        RECT 117.585 195.625 118.045 196.675 ;
        RECT 115.860 195.315 116.715 195.485 ;
        RECT 116.920 195.315 117.415 195.485 ;
        RECT 117.585 195.095 117.915 195.455 ;
        RECT 118.275 195.355 118.445 197.475 ;
        RECT 118.615 197.145 118.945 197.645 ;
        RECT 119.115 196.975 119.370 197.475 ;
        RECT 118.620 196.805 119.370 196.975 ;
        RECT 118.620 195.815 118.850 196.805 ;
        RECT 119.020 195.985 119.370 196.635 ;
        RECT 119.545 196.555 120.755 197.645 ;
        RECT 120.930 197.210 126.275 197.645 ;
        RECT 119.545 196.015 120.065 196.555 ;
        RECT 120.235 195.845 120.755 196.385 ;
        RECT 122.520 195.960 122.870 197.210 ;
        RECT 126.445 196.555 127.655 197.645 ;
        RECT 118.620 195.645 119.370 195.815 ;
        RECT 118.615 195.095 118.945 195.475 ;
        RECT 119.115 195.355 119.370 195.645 ;
        RECT 119.545 195.095 120.755 195.845 ;
        RECT 124.350 195.640 124.690 196.470 ;
        RECT 126.445 196.015 126.965 196.555 ;
        RECT 127.135 195.845 127.655 196.385 ;
        RECT 120.930 195.095 126.275 195.640 ;
        RECT 126.445 195.095 127.655 195.845 ;
        RECT 14.580 194.925 127.740 195.095 ;
        RECT 14.665 194.175 15.875 194.925 ;
        RECT 14.665 193.635 15.185 194.175 ;
        RECT 16.965 194.155 20.475 194.925 ;
        RECT 20.650 194.380 25.995 194.925 ;
        RECT 26.170 194.380 31.515 194.925 ;
        RECT 31.690 194.380 37.035 194.925 ;
        RECT 15.355 193.465 15.875 194.005 ;
        RECT 14.665 192.375 15.875 193.465 ;
        RECT 16.965 193.465 18.655 193.985 ;
        RECT 18.825 193.635 20.475 194.155 ;
        RECT 16.965 192.375 20.475 193.465 ;
        RECT 22.240 192.810 22.590 194.060 ;
        RECT 24.070 193.550 24.410 194.380 ;
        RECT 27.760 192.810 28.110 194.060 ;
        RECT 29.590 193.550 29.930 194.380 ;
        RECT 33.280 192.810 33.630 194.060 ;
        RECT 35.110 193.550 35.450 194.380 ;
        RECT 37.205 194.200 37.495 194.925 ;
        RECT 38.585 194.155 42.095 194.925 ;
        RECT 42.270 194.380 47.615 194.925 ;
        RECT 20.650 192.375 25.995 192.810 ;
        RECT 26.170 192.375 31.515 192.810 ;
        RECT 31.690 192.375 37.035 192.810 ;
        RECT 37.205 192.375 37.495 193.540 ;
        RECT 38.585 193.465 40.275 193.985 ;
        RECT 40.445 193.635 42.095 194.155 ;
        RECT 38.585 192.375 42.095 193.465 ;
        RECT 43.860 192.810 44.210 194.060 ;
        RECT 45.690 193.550 46.030 194.380 ;
        RECT 47.845 194.105 48.055 194.925 ;
        RECT 48.225 194.125 48.555 194.755 ;
        RECT 48.225 193.525 48.475 194.125 ;
        RECT 48.725 194.105 48.955 194.925 ;
        RECT 49.170 194.375 49.425 194.665 ;
        RECT 49.595 194.545 49.925 194.925 ;
        RECT 49.170 194.205 49.920 194.375 ;
        RECT 48.645 193.685 48.975 193.935 ;
        RECT 42.270 192.375 47.615 192.810 ;
        RECT 47.845 192.375 48.055 193.515 ;
        RECT 48.225 192.545 48.555 193.525 ;
        RECT 48.725 192.375 48.955 193.515 ;
        RECT 49.170 193.385 49.520 194.035 ;
        RECT 49.690 193.215 49.920 194.205 ;
        RECT 49.170 193.045 49.920 193.215 ;
        RECT 49.170 192.545 49.425 193.045 ;
        RECT 49.595 192.375 49.925 192.875 ;
        RECT 50.095 192.545 50.265 194.665 ;
        RECT 50.625 194.565 50.955 194.925 ;
        RECT 51.125 194.535 51.620 194.705 ;
        RECT 51.825 194.535 52.680 194.705 ;
        RECT 50.495 193.345 50.955 194.395 ;
        RECT 50.435 192.560 50.760 193.345 ;
        RECT 51.125 193.175 51.295 194.535 ;
        RECT 51.465 193.625 51.815 194.245 ;
        RECT 51.985 194.025 52.340 194.245 ;
        RECT 51.985 193.435 52.155 194.025 ;
        RECT 52.510 193.825 52.680 194.535 ;
        RECT 53.555 194.465 53.885 194.925 ;
        RECT 54.095 194.565 54.445 194.735 ;
        RECT 52.885 193.995 53.675 194.245 ;
        RECT 54.095 194.175 54.355 194.565 ;
        RECT 54.665 194.475 55.615 194.755 ;
        RECT 55.785 194.485 55.975 194.925 ;
        RECT 56.145 194.545 57.215 194.715 ;
        RECT 53.845 193.825 54.015 194.005 ;
        RECT 51.125 193.005 51.520 193.175 ;
        RECT 51.690 193.045 52.155 193.435 ;
        RECT 52.325 193.655 54.015 193.825 ;
        RECT 51.350 192.875 51.520 193.005 ;
        RECT 52.325 192.875 52.495 193.655 ;
        RECT 54.185 193.485 54.355 194.175 ;
        RECT 52.855 193.315 54.355 193.485 ;
        RECT 54.545 193.515 54.755 194.305 ;
        RECT 54.925 193.685 55.275 194.305 ;
        RECT 55.445 193.695 55.615 194.475 ;
        RECT 56.145 194.315 56.315 194.545 ;
        RECT 55.785 194.145 56.315 194.315 ;
        RECT 55.785 193.865 56.005 194.145 ;
        RECT 56.485 193.975 56.725 194.375 ;
        RECT 55.445 193.525 55.850 193.695 ;
        RECT 56.185 193.605 56.725 193.975 ;
        RECT 56.895 194.190 57.215 194.545 ;
        RECT 57.460 194.465 57.765 194.925 ;
        RECT 57.935 194.215 58.190 194.745 ;
        RECT 56.895 194.015 57.220 194.190 ;
        RECT 56.895 193.715 57.810 194.015 ;
        RECT 57.070 193.685 57.810 193.715 ;
        RECT 54.545 193.355 55.220 193.515 ;
        RECT 55.680 193.435 55.850 193.525 ;
        RECT 54.545 193.345 55.510 193.355 ;
        RECT 54.185 193.175 54.355 193.315 ;
        RECT 50.930 192.375 51.180 192.835 ;
        RECT 51.350 192.545 51.600 192.875 ;
        RECT 51.815 192.545 52.495 192.875 ;
        RECT 52.665 192.975 53.740 193.145 ;
        RECT 54.185 193.005 54.745 193.175 ;
        RECT 55.050 193.055 55.510 193.345 ;
        RECT 55.680 193.265 56.900 193.435 ;
        RECT 52.665 192.635 52.835 192.975 ;
        RECT 53.070 192.375 53.400 192.805 ;
        RECT 53.570 192.635 53.740 192.975 ;
        RECT 54.035 192.375 54.405 192.835 ;
        RECT 54.575 192.545 54.745 193.005 ;
        RECT 55.680 192.885 55.850 193.265 ;
        RECT 57.070 193.095 57.240 193.685 ;
        RECT 57.980 193.565 58.190 194.215 ;
        RECT 59.285 194.155 62.795 194.925 ;
        RECT 62.965 194.200 63.255 194.925 ;
        RECT 63.425 194.155 65.095 194.925 ;
        RECT 54.980 192.545 55.850 192.885 ;
        RECT 56.440 192.925 57.240 193.095 ;
        RECT 56.020 192.375 56.270 192.835 ;
        RECT 56.440 192.635 56.610 192.925 ;
        RECT 56.790 192.375 57.120 192.755 ;
        RECT 57.460 192.375 57.765 193.515 ;
        RECT 57.935 192.685 58.190 193.565 ;
        RECT 59.285 193.465 60.975 193.985 ;
        RECT 61.145 193.635 62.795 194.155 ;
        RECT 59.285 192.375 62.795 193.465 ;
        RECT 62.965 192.375 63.255 193.540 ;
        RECT 63.425 193.465 64.175 193.985 ;
        RECT 64.345 193.635 65.095 194.155 ;
        RECT 65.325 194.105 65.535 194.925 ;
        RECT 65.705 194.125 66.035 194.755 ;
        RECT 65.705 193.525 65.955 194.125 ;
        RECT 66.205 194.105 66.435 194.925 ;
        RECT 67.105 194.155 68.775 194.925 ;
        RECT 66.125 193.685 66.455 193.935 ;
        RECT 63.425 192.375 65.095 193.465 ;
        RECT 65.325 192.375 65.535 193.515 ;
        RECT 65.705 192.545 66.035 193.525 ;
        RECT 66.205 192.375 66.435 193.515 ;
        RECT 67.105 193.465 67.855 193.985 ;
        RECT 68.025 193.635 68.775 194.155 ;
        RECT 68.945 194.105 69.205 194.925 ;
        RECT 69.375 194.105 69.705 194.525 ;
        RECT 69.885 194.355 70.145 194.755 ;
        RECT 70.315 194.525 70.645 194.925 ;
        RECT 70.815 194.355 70.985 194.705 ;
        RECT 71.155 194.525 71.530 194.925 ;
        RECT 69.885 194.185 71.550 194.355 ;
        RECT 71.720 194.250 71.995 194.595 ;
        RECT 69.455 194.015 69.705 194.105 ;
        RECT 71.380 194.015 71.550 194.185 ;
        RECT 68.950 193.685 69.285 193.935 ;
        RECT 69.455 193.685 70.170 194.015 ;
        RECT 70.385 193.685 71.210 194.015 ;
        RECT 71.380 193.685 71.655 194.015 ;
        RECT 67.105 192.375 68.775 193.465 ;
        RECT 68.945 192.375 69.205 193.515 ;
        RECT 69.455 193.125 69.625 193.685 ;
        RECT 69.885 193.225 70.215 193.515 ;
        RECT 70.385 193.395 70.630 193.685 ;
        RECT 71.380 193.515 71.550 193.685 ;
        RECT 71.825 193.515 71.995 194.250 ;
        RECT 70.890 193.345 71.550 193.515 ;
        RECT 70.890 193.225 71.060 193.345 ;
        RECT 69.885 193.055 71.060 193.225 ;
        RECT 69.445 192.555 71.060 192.885 ;
        RECT 71.230 192.375 71.510 193.175 ;
        RECT 71.720 192.545 71.995 193.515 ;
        RECT 72.165 194.250 72.440 194.595 ;
        RECT 72.630 194.525 73.005 194.925 ;
        RECT 73.175 194.355 73.345 194.705 ;
        RECT 73.515 194.525 73.845 194.925 ;
        RECT 74.015 194.355 74.275 194.755 ;
        RECT 72.165 193.515 72.335 194.250 ;
        RECT 72.610 194.185 74.275 194.355 ;
        RECT 72.610 194.015 72.780 194.185 ;
        RECT 74.455 194.105 74.785 194.525 ;
        RECT 74.955 194.105 75.215 194.925 ;
        RECT 75.385 194.155 78.895 194.925 ;
        RECT 79.070 194.380 84.415 194.925 ;
        RECT 74.455 194.015 74.705 194.105 ;
        RECT 72.505 193.685 72.780 194.015 ;
        RECT 72.950 193.685 73.775 194.015 ;
        RECT 73.990 193.685 74.705 194.015 ;
        RECT 74.875 193.685 75.210 193.935 ;
        RECT 72.610 193.515 72.780 193.685 ;
        RECT 72.165 192.545 72.440 193.515 ;
        RECT 72.610 193.345 73.270 193.515 ;
        RECT 73.530 193.395 73.775 193.685 ;
        RECT 73.100 193.225 73.270 193.345 ;
        RECT 73.945 193.225 74.275 193.515 ;
        RECT 72.650 192.375 72.930 193.175 ;
        RECT 73.100 193.055 74.275 193.225 ;
        RECT 74.535 193.125 74.705 193.685 ;
        RECT 73.100 192.555 74.715 192.885 ;
        RECT 74.955 192.375 75.215 193.515 ;
        RECT 75.385 193.465 77.075 193.985 ;
        RECT 77.245 193.635 78.895 194.155 ;
        RECT 75.385 192.375 78.895 193.465 ;
        RECT 80.660 192.810 81.010 194.060 ;
        RECT 82.490 193.550 82.830 194.380 ;
        RECT 84.860 194.115 85.105 194.720 ;
        RECT 85.325 194.390 85.835 194.925 ;
        RECT 84.585 193.945 85.815 194.115 ;
        RECT 84.585 193.135 84.925 193.945 ;
        RECT 85.095 193.380 85.845 193.570 ;
        RECT 79.070 192.375 84.415 192.810 ;
        RECT 84.585 192.725 85.100 193.135 ;
        RECT 85.335 192.375 85.505 193.135 ;
        RECT 85.675 192.715 85.845 193.380 ;
        RECT 86.015 193.395 86.205 194.755 ;
        RECT 86.375 193.905 86.650 194.755 ;
        RECT 86.840 194.390 87.370 194.755 ;
        RECT 87.795 194.525 88.125 194.925 ;
        RECT 87.195 194.355 87.370 194.390 ;
        RECT 86.375 193.735 86.655 193.905 ;
        RECT 86.375 193.595 86.650 193.735 ;
        RECT 86.855 193.395 87.025 194.195 ;
        RECT 86.015 193.225 87.025 193.395 ;
        RECT 87.195 194.185 88.125 194.355 ;
        RECT 88.295 194.185 88.550 194.755 ;
        RECT 88.725 194.200 89.015 194.925 ;
        RECT 87.195 193.055 87.365 194.185 ;
        RECT 87.955 194.015 88.125 194.185 ;
        RECT 86.240 192.885 87.365 193.055 ;
        RECT 87.535 193.685 87.730 194.015 ;
        RECT 87.955 193.685 88.210 194.015 ;
        RECT 87.535 192.715 87.705 193.685 ;
        RECT 88.380 193.515 88.550 194.185 ;
        RECT 89.245 194.105 89.455 194.925 ;
        RECT 89.625 194.125 89.955 194.755 ;
        RECT 85.675 192.545 87.705 192.715 ;
        RECT 87.875 192.375 88.045 193.515 ;
        RECT 88.215 192.545 88.550 193.515 ;
        RECT 88.725 192.375 89.015 193.540 ;
        RECT 89.625 193.525 89.875 194.125 ;
        RECT 90.125 194.105 90.355 194.925 ;
        RECT 90.565 194.155 93.155 194.925 ;
        RECT 90.045 193.685 90.375 193.935 ;
        RECT 89.245 192.375 89.455 193.515 ;
        RECT 89.625 192.545 89.955 193.525 ;
        RECT 90.125 192.375 90.355 193.515 ;
        RECT 90.565 193.465 91.775 193.985 ;
        RECT 91.945 193.635 93.155 194.155 ;
        RECT 93.365 194.105 93.595 194.925 ;
        RECT 93.765 194.125 94.095 194.755 ;
        RECT 93.345 193.685 93.675 193.935 ;
        RECT 93.845 193.525 94.095 194.125 ;
        RECT 94.265 194.105 94.475 194.925 ;
        RECT 94.705 194.415 95.010 194.925 ;
        RECT 94.705 193.685 95.020 194.245 ;
        RECT 95.190 193.935 95.440 194.745 ;
        RECT 95.610 194.400 95.870 194.925 ;
        RECT 96.050 193.935 96.300 194.745 ;
        RECT 96.470 194.365 96.730 194.925 ;
        RECT 96.900 194.275 97.160 194.730 ;
        RECT 97.330 194.445 97.590 194.925 ;
        RECT 97.760 194.275 98.020 194.730 ;
        RECT 98.190 194.445 98.450 194.925 ;
        RECT 98.620 194.275 98.880 194.730 ;
        RECT 99.050 194.445 99.295 194.925 ;
        RECT 99.465 194.275 99.740 194.730 ;
        RECT 99.910 194.445 100.155 194.925 ;
        RECT 100.325 194.275 100.585 194.730 ;
        RECT 100.765 194.445 101.015 194.925 ;
        RECT 101.185 194.275 101.445 194.730 ;
        RECT 101.625 194.445 101.875 194.925 ;
        RECT 102.045 194.275 102.305 194.730 ;
        RECT 102.485 194.445 102.745 194.925 ;
        RECT 102.915 194.275 103.175 194.730 ;
        RECT 103.345 194.445 103.645 194.925 ;
        RECT 96.900 194.245 103.645 194.275 ;
        RECT 96.900 194.105 103.675 194.245 ;
        RECT 103.905 194.175 105.115 194.925 ;
        RECT 102.480 194.075 103.675 194.105 ;
        RECT 95.190 193.685 102.310 193.935 ;
        RECT 90.565 192.375 93.155 193.465 ;
        RECT 93.365 192.375 93.595 193.515 ;
        RECT 93.765 192.545 94.095 193.525 ;
        RECT 94.265 192.375 94.475 193.515 ;
        RECT 94.715 192.375 95.010 193.185 ;
        RECT 95.190 192.545 95.435 193.685 ;
        RECT 95.610 192.375 95.870 193.185 ;
        RECT 96.050 192.550 96.300 193.685 ;
        RECT 102.480 193.515 103.645 194.075 ;
        RECT 96.900 193.290 103.645 193.515 ;
        RECT 103.905 193.465 104.425 194.005 ;
        RECT 104.595 193.635 105.115 194.175 ;
        RECT 105.285 194.155 108.795 194.925 ;
        RECT 105.285 193.465 106.975 193.985 ;
        RECT 107.145 193.635 108.795 194.155 ;
        RECT 109.005 194.105 109.235 194.925 ;
        RECT 109.405 194.125 109.735 194.755 ;
        RECT 108.985 193.685 109.315 193.935 ;
        RECT 109.485 193.525 109.735 194.125 ;
        RECT 109.905 194.105 110.115 194.925 ;
        RECT 110.620 194.115 110.865 194.720 ;
        RECT 111.085 194.390 111.595 194.925 ;
        RECT 96.900 193.275 102.305 193.290 ;
        RECT 96.470 192.380 96.730 193.175 ;
        RECT 96.900 192.550 97.160 193.275 ;
        RECT 97.330 192.380 97.590 193.105 ;
        RECT 97.760 192.550 98.020 193.275 ;
        RECT 98.190 192.380 98.450 193.105 ;
        RECT 98.620 192.550 98.880 193.275 ;
        RECT 99.050 192.380 99.310 193.105 ;
        RECT 99.480 192.550 99.740 193.275 ;
        RECT 99.910 192.380 100.155 193.105 ;
        RECT 100.325 192.550 100.585 193.275 ;
        RECT 100.770 192.380 101.015 193.105 ;
        RECT 101.185 192.550 101.445 193.275 ;
        RECT 101.630 192.380 101.875 193.105 ;
        RECT 102.045 192.550 102.305 193.275 ;
        RECT 102.490 192.380 102.745 193.105 ;
        RECT 102.915 192.550 103.205 193.290 ;
        RECT 96.470 192.375 102.745 192.380 ;
        RECT 103.375 192.375 103.645 193.120 ;
        RECT 103.905 192.375 105.115 193.465 ;
        RECT 105.285 192.375 108.795 193.465 ;
        RECT 109.005 192.375 109.235 193.515 ;
        RECT 109.405 192.545 109.735 193.525 ;
        RECT 110.345 193.945 111.575 194.115 ;
        RECT 109.905 192.375 110.115 193.515 ;
        RECT 110.345 193.135 110.685 193.945 ;
        RECT 110.855 193.380 111.605 193.570 ;
        RECT 110.345 192.725 110.860 193.135 ;
        RECT 111.095 192.375 111.265 193.135 ;
        RECT 111.435 192.715 111.605 193.380 ;
        RECT 111.775 193.395 111.965 194.755 ;
        RECT 112.135 194.585 112.410 194.755 ;
        RECT 112.135 194.415 112.415 194.585 ;
        RECT 112.135 193.595 112.410 194.415 ;
        RECT 112.600 194.390 113.130 194.755 ;
        RECT 113.555 194.525 113.885 194.925 ;
        RECT 112.955 194.355 113.130 194.390 ;
        RECT 112.615 193.395 112.785 194.195 ;
        RECT 111.775 193.225 112.785 193.395 ;
        RECT 112.955 194.185 113.885 194.355 ;
        RECT 114.055 194.185 114.310 194.755 ;
        RECT 114.485 194.200 114.775 194.925 ;
        RECT 112.955 193.055 113.125 194.185 ;
        RECT 113.715 194.015 113.885 194.185 ;
        RECT 112.000 192.885 113.125 193.055 ;
        RECT 113.295 193.685 113.490 194.015 ;
        RECT 113.715 193.685 113.970 194.015 ;
        RECT 113.295 192.715 113.465 193.685 ;
        RECT 114.140 193.515 114.310 194.185 ;
        RECT 115.005 194.105 115.215 194.925 ;
        RECT 115.385 194.125 115.715 194.755 ;
        RECT 111.435 192.545 113.465 192.715 ;
        RECT 113.635 192.375 113.805 193.515 ;
        RECT 113.975 192.545 114.310 193.515 ;
        RECT 114.485 192.375 114.775 193.540 ;
        RECT 115.385 193.525 115.635 194.125 ;
        RECT 115.885 194.105 116.115 194.925 ;
        RECT 117.245 194.155 120.755 194.925 ;
        RECT 120.930 194.380 126.275 194.925 ;
        RECT 115.805 193.685 116.135 193.935 ;
        RECT 115.005 192.375 115.215 193.515 ;
        RECT 115.385 192.545 115.715 193.525 ;
        RECT 115.885 192.375 116.115 193.515 ;
        RECT 117.245 193.465 118.935 193.985 ;
        RECT 119.105 193.635 120.755 194.155 ;
        RECT 117.245 192.375 120.755 193.465 ;
        RECT 122.520 192.810 122.870 194.060 ;
        RECT 124.350 193.550 124.690 194.380 ;
        RECT 126.445 194.175 127.655 194.925 ;
        RECT 126.445 193.465 126.965 194.005 ;
        RECT 127.135 193.635 127.655 194.175 ;
        RECT 120.930 192.375 126.275 192.810 ;
        RECT 126.445 192.375 127.655 193.465 ;
        RECT 14.580 192.205 127.740 192.375 ;
        RECT 14.665 191.115 15.875 192.205 ;
        RECT 14.665 190.405 15.185 190.945 ;
        RECT 15.355 190.575 15.875 191.115 ;
        RECT 16.045 191.115 18.635 192.205 ;
        RECT 18.810 191.770 24.155 192.205 ;
        RECT 16.045 190.595 17.255 191.115 ;
        RECT 17.425 190.425 18.635 190.945 ;
        RECT 20.400 190.520 20.750 191.770 ;
        RECT 24.325 191.040 24.615 192.205 ;
        RECT 25.250 191.770 30.595 192.205 ;
        RECT 30.770 191.770 36.115 192.205 ;
        RECT 14.665 189.655 15.875 190.405 ;
        RECT 16.045 189.655 18.635 190.425 ;
        RECT 22.230 190.200 22.570 191.030 ;
        RECT 26.840 190.520 27.190 191.770 ;
        RECT 18.810 189.655 24.155 190.200 ;
        RECT 24.325 189.655 24.615 190.380 ;
        RECT 28.670 190.200 29.010 191.030 ;
        RECT 32.360 190.520 32.710 191.770 ;
        RECT 36.660 191.225 36.915 191.895 ;
        RECT 37.095 191.405 37.380 192.205 ;
        RECT 37.560 191.485 37.890 191.995 ;
        RECT 36.660 191.185 36.840 191.225 ;
        RECT 34.190 190.200 34.530 191.030 ;
        RECT 36.575 191.015 36.840 191.185 ;
        RECT 36.660 190.365 36.840 191.015 ;
        RECT 37.560 190.895 37.810 191.485 ;
        RECT 38.160 191.335 38.330 191.945 ;
        RECT 38.500 191.515 38.830 192.205 ;
        RECT 39.060 191.655 39.300 191.945 ;
        RECT 39.500 191.825 39.920 192.205 ;
        RECT 40.100 191.735 40.730 191.985 ;
        RECT 41.200 191.825 41.530 192.205 ;
        RECT 40.100 191.655 40.270 191.735 ;
        RECT 41.700 191.655 41.870 191.945 ;
        RECT 42.050 191.825 42.430 192.205 ;
        RECT 42.670 191.820 43.500 191.990 ;
        RECT 39.060 191.485 40.270 191.655 ;
        RECT 37.010 190.565 37.810 190.895 ;
        RECT 25.250 189.655 30.595 190.200 ;
        RECT 30.770 189.655 36.115 190.200 ;
        RECT 36.660 189.835 36.915 190.365 ;
        RECT 37.095 189.655 37.380 190.115 ;
        RECT 37.560 189.915 37.810 190.565 ;
        RECT 38.010 191.315 38.330 191.335 ;
        RECT 38.010 191.145 39.930 191.315 ;
        RECT 38.010 190.250 38.200 191.145 ;
        RECT 40.100 190.975 40.270 191.485 ;
        RECT 40.440 191.225 40.960 191.535 ;
        RECT 38.370 190.805 40.270 190.975 ;
        RECT 38.370 190.745 38.700 190.805 ;
        RECT 38.850 190.575 39.180 190.635 ;
        RECT 38.520 190.305 39.180 190.575 ;
        RECT 38.010 189.920 38.330 190.250 ;
        RECT 38.510 189.655 39.170 190.135 ;
        RECT 39.370 190.045 39.540 190.805 ;
        RECT 40.440 190.635 40.620 191.045 ;
        RECT 39.710 190.465 40.040 190.585 ;
        RECT 40.790 190.465 40.960 191.225 ;
        RECT 39.710 190.295 40.960 190.465 ;
        RECT 41.130 191.405 42.500 191.655 ;
        RECT 41.130 190.635 41.320 191.405 ;
        RECT 42.250 191.145 42.500 191.405 ;
        RECT 41.490 190.975 41.740 191.135 ;
        RECT 42.670 190.975 42.840 191.820 ;
        RECT 43.735 191.535 43.905 192.035 ;
        RECT 44.075 191.705 44.405 192.205 ;
        RECT 43.010 191.145 43.510 191.525 ;
        RECT 43.735 191.365 44.430 191.535 ;
        RECT 41.490 190.805 42.840 190.975 ;
        RECT 42.420 190.765 42.840 190.805 ;
        RECT 41.130 190.295 41.550 190.635 ;
        RECT 41.840 190.305 42.250 190.635 ;
        RECT 39.370 189.875 40.220 190.045 ;
        RECT 40.780 189.655 41.100 190.115 ;
        RECT 41.300 189.865 41.550 190.295 ;
        RECT 41.840 189.655 42.250 190.095 ;
        RECT 42.420 190.035 42.590 190.765 ;
        RECT 42.760 190.215 43.110 190.585 ;
        RECT 43.290 190.275 43.510 191.145 ;
        RECT 43.680 190.575 44.090 191.195 ;
        RECT 44.260 190.395 44.430 191.365 ;
        RECT 43.735 190.205 44.430 190.395 ;
        RECT 42.420 189.835 43.435 190.035 ;
        RECT 43.735 189.875 43.905 190.205 ;
        RECT 44.075 189.655 44.405 190.035 ;
        RECT 44.620 189.915 44.845 192.035 ;
        RECT 45.015 191.705 45.345 192.205 ;
        RECT 45.515 191.535 45.685 192.035 ;
        RECT 45.020 191.365 45.685 191.535 ;
        RECT 45.945 191.445 46.460 191.855 ;
        RECT 46.695 191.445 46.865 192.205 ;
        RECT 47.035 191.865 49.065 192.035 ;
        RECT 45.020 190.375 45.250 191.365 ;
        RECT 45.420 190.545 45.770 191.195 ;
        RECT 45.945 190.635 46.285 191.445 ;
        RECT 47.035 191.200 47.205 191.865 ;
        RECT 47.600 191.525 48.725 191.695 ;
        RECT 46.455 191.010 47.205 191.200 ;
        RECT 47.375 191.185 48.385 191.355 ;
        RECT 45.945 190.465 47.175 190.635 ;
        RECT 45.020 190.205 45.685 190.375 ;
        RECT 45.015 189.655 45.345 190.035 ;
        RECT 45.515 189.915 45.685 190.205 ;
        RECT 46.220 189.860 46.465 190.465 ;
        RECT 46.685 189.655 47.195 190.190 ;
        RECT 47.375 189.825 47.565 191.185 ;
        RECT 47.735 190.845 48.010 190.985 ;
        RECT 47.735 190.675 48.015 190.845 ;
        RECT 47.735 189.825 48.010 190.675 ;
        RECT 48.215 190.385 48.385 191.185 ;
        RECT 48.555 190.395 48.725 191.525 ;
        RECT 48.895 190.895 49.065 191.865 ;
        RECT 49.235 191.065 49.405 192.205 ;
        RECT 49.575 191.065 49.910 192.035 ;
        RECT 48.895 190.565 49.090 190.895 ;
        RECT 49.315 190.565 49.570 190.895 ;
        RECT 49.315 190.395 49.485 190.565 ;
        RECT 49.740 190.395 49.910 191.065 ;
        RECT 50.085 191.040 50.375 192.205 ;
        RECT 51.005 191.130 51.275 192.035 ;
        RECT 51.445 191.445 51.775 192.205 ;
        RECT 51.955 191.275 52.125 192.035 ;
        RECT 48.555 190.225 49.485 190.395 ;
        RECT 48.555 190.190 48.730 190.225 ;
        RECT 48.200 189.825 48.730 190.190 ;
        RECT 49.155 189.655 49.485 190.055 ;
        RECT 49.655 189.825 49.910 190.395 ;
        RECT 50.085 189.655 50.375 190.380 ;
        RECT 51.005 190.330 51.175 191.130 ;
        RECT 51.460 191.105 52.125 191.275 ;
        RECT 51.460 190.960 51.630 191.105 ;
        RECT 51.345 190.630 51.630 190.960 ;
        RECT 52.390 191.015 52.645 191.895 ;
        RECT 52.815 191.065 53.120 192.205 ;
        RECT 53.460 191.825 53.790 192.205 ;
        RECT 53.970 191.655 54.140 191.945 ;
        RECT 54.310 191.745 54.560 192.205 ;
        RECT 53.340 191.485 54.140 191.655 ;
        RECT 54.730 191.695 55.600 192.035 ;
        RECT 51.460 190.375 51.630 190.630 ;
        RECT 51.865 190.555 52.195 190.925 ;
        RECT 51.005 189.825 51.265 190.330 ;
        RECT 51.460 190.205 52.125 190.375 ;
        RECT 51.445 189.655 51.775 190.035 ;
        RECT 51.955 189.825 52.125 190.205 ;
        RECT 52.390 190.365 52.600 191.015 ;
        RECT 53.340 190.895 53.510 191.485 ;
        RECT 54.730 191.315 54.900 191.695 ;
        RECT 55.835 191.575 56.005 192.035 ;
        RECT 56.175 191.745 56.545 192.205 ;
        RECT 56.840 191.605 57.010 191.945 ;
        RECT 57.180 191.775 57.510 192.205 ;
        RECT 57.745 191.605 57.915 191.945 ;
        RECT 53.680 191.145 54.900 191.315 ;
        RECT 55.070 191.235 55.530 191.525 ;
        RECT 55.835 191.405 56.395 191.575 ;
        RECT 56.840 191.435 57.915 191.605 ;
        RECT 58.085 191.705 58.765 192.035 ;
        RECT 58.980 191.705 59.230 192.035 ;
        RECT 59.400 191.745 59.650 192.205 ;
        RECT 56.225 191.265 56.395 191.405 ;
        RECT 55.070 191.225 56.035 191.235 ;
        RECT 54.730 191.055 54.900 191.145 ;
        RECT 55.360 191.065 56.035 191.225 ;
        RECT 52.770 190.865 53.510 190.895 ;
        RECT 52.770 190.565 53.685 190.865 ;
        RECT 53.360 190.390 53.685 190.565 ;
        RECT 52.390 189.835 52.645 190.365 ;
        RECT 52.815 189.655 53.120 190.115 ;
        RECT 53.365 190.035 53.685 190.390 ;
        RECT 53.855 190.605 54.395 190.975 ;
        RECT 54.730 190.885 55.135 191.055 ;
        RECT 53.855 190.205 54.095 190.605 ;
        RECT 54.575 190.435 54.795 190.715 ;
        RECT 54.265 190.265 54.795 190.435 ;
        RECT 54.265 190.035 54.435 190.265 ;
        RECT 54.965 190.105 55.135 190.885 ;
        RECT 55.305 190.275 55.655 190.895 ;
        RECT 55.825 190.275 56.035 191.065 ;
        RECT 56.225 191.095 57.725 191.265 ;
        RECT 56.225 190.405 56.395 191.095 ;
        RECT 58.085 190.925 58.255 191.705 ;
        RECT 59.060 191.575 59.230 191.705 ;
        RECT 56.565 190.755 58.255 190.925 ;
        RECT 58.425 191.145 58.890 191.535 ;
        RECT 59.060 191.405 59.455 191.575 ;
        RECT 56.565 190.575 56.735 190.755 ;
        RECT 53.365 189.865 54.435 190.035 ;
        RECT 54.605 189.655 54.795 190.095 ;
        RECT 54.965 189.825 55.915 190.105 ;
        RECT 56.225 190.015 56.485 190.405 ;
        RECT 56.905 190.335 57.695 190.585 ;
        RECT 56.135 189.845 56.485 190.015 ;
        RECT 56.695 189.655 57.025 190.115 ;
        RECT 57.900 190.045 58.070 190.755 ;
        RECT 58.425 190.555 58.595 191.145 ;
        RECT 58.240 190.335 58.595 190.555 ;
        RECT 58.765 190.335 59.115 190.955 ;
        RECT 59.285 190.045 59.455 191.405 ;
        RECT 59.820 191.235 60.145 192.020 ;
        RECT 59.625 190.185 60.085 191.235 ;
        RECT 57.900 189.875 58.755 190.045 ;
        RECT 58.960 189.875 59.455 190.045 ;
        RECT 59.625 189.655 59.955 190.015 ;
        RECT 60.315 189.915 60.485 192.035 ;
        RECT 60.655 191.705 60.985 192.205 ;
        RECT 61.155 191.535 61.410 192.035 ;
        RECT 60.660 191.365 61.410 191.535 ;
        RECT 60.660 190.375 60.890 191.365 ;
        RECT 61.060 190.545 61.410 191.195 ;
        RECT 61.635 191.065 61.885 192.205 ;
        RECT 62.055 191.015 62.305 191.895 ;
        RECT 62.475 191.065 62.780 192.205 ;
        RECT 63.120 191.825 63.450 192.205 ;
        RECT 63.630 191.655 63.800 191.945 ;
        RECT 63.970 191.745 64.220 192.205 ;
        RECT 63.000 191.485 63.800 191.655 ;
        RECT 64.390 191.695 65.260 192.035 ;
        RECT 60.660 190.205 61.410 190.375 ;
        RECT 60.655 189.655 60.985 190.035 ;
        RECT 61.155 189.915 61.410 190.205 ;
        RECT 61.635 189.655 61.885 190.410 ;
        RECT 62.055 190.365 62.260 191.015 ;
        RECT 63.000 190.895 63.170 191.485 ;
        RECT 64.390 191.315 64.560 191.695 ;
        RECT 65.495 191.575 65.665 192.035 ;
        RECT 65.835 191.745 66.205 192.205 ;
        RECT 66.500 191.605 66.670 191.945 ;
        RECT 66.840 191.775 67.170 192.205 ;
        RECT 67.405 191.605 67.575 191.945 ;
        RECT 63.340 191.145 64.560 191.315 ;
        RECT 64.730 191.235 65.190 191.525 ;
        RECT 65.495 191.405 66.055 191.575 ;
        RECT 66.500 191.435 67.575 191.605 ;
        RECT 67.745 191.705 68.425 192.035 ;
        RECT 68.640 191.705 68.890 192.035 ;
        RECT 69.060 191.745 69.310 192.205 ;
        RECT 65.885 191.265 66.055 191.405 ;
        RECT 64.730 191.225 65.695 191.235 ;
        RECT 64.390 191.055 64.560 191.145 ;
        RECT 65.020 191.065 65.695 191.225 ;
        RECT 62.430 190.865 63.170 190.895 ;
        RECT 62.430 190.565 63.345 190.865 ;
        RECT 63.020 190.390 63.345 190.565 ;
        RECT 62.055 189.835 62.305 190.365 ;
        RECT 62.475 189.655 62.780 190.115 ;
        RECT 63.025 190.035 63.345 190.390 ;
        RECT 63.515 190.605 64.055 190.975 ;
        RECT 64.390 190.885 64.795 191.055 ;
        RECT 63.515 190.205 63.755 190.605 ;
        RECT 64.235 190.435 64.455 190.715 ;
        RECT 63.925 190.265 64.455 190.435 ;
        RECT 63.925 190.035 64.095 190.265 ;
        RECT 64.625 190.105 64.795 190.885 ;
        RECT 64.965 190.275 65.315 190.895 ;
        RECT 65.485 190.275 65.695 191.065 ;
        RECT 65.885 191.095 67.385 191.265 ;
        RECT 65.885 190.405 66.055 191.095 ;
        RECT 67.745 190.925 67.915 191.705 ;
        RECT 68.720 191.575 68.890 191.705 ;
        RECT 66.225 190.755 67.915 190.925 ;
        RECT 68.085 191.145 68.550 191.535 ;
        RECT 68.720 191.405 69.115 191.575 ;
        RECT 66.225 190.575 66.395 190.755 ;
        RECT 63.025 189.865 64.095 190.035 ;
        RECT 64.265 189.655 64.455 190.095 ;
        RECT 64.625 189.825 65.575 190.105 ;
        RECT 65.885 190.015 66.145 190.405 ;
        RECT 66.565 190.335 67.355 190.585 ;
        RECT 65.795 189.845 66.145 190.015 ;
        RECT 66.355 189.655 66.685 190.115 ;
        RECT 67.560 190.045 67.730 190.755 ;
        RECT 68.085 190.555 68.255 191.145 ;
        RECT 67.900 190.335 68.255 190.555 ;
        RECT 68.425 190.335 68.775 190.955 ;
        RECT 68.945 190.045 69.115 191.405 ;
        RECT 69.480 191.235 69.805 192.020 ;
        RECT 69.285 190.185 69.745 191.235 ;
        RECT 67.560 189.875 68.415 190.045 ;
        RECT 68.620 189.875 69.115 190.045 ;
        RECT 69.285 189.655 69.615 190.015 ;
        RECT 69.975 189.915 70.145 192.035 ;
        RECT 70.315 191.705 70.645 192.205 ;
        RECT 70.815 191.535 71.070 192.035 ;
        RECT 71.265 191.695 71.565 192.205 ;
        RECT 71.735 191.695 72.115 191.865 ;
        RECT 72.695 191.695 73.325 192.205 ;
        RECT 70.320 191.365 71.070 191.535 ;
        RECT 71.735 191.525 71.905 191.695 ;
        RECT 73.495 191.525 73.825 192.035 ;
        RECT 73.995 191.695 74.295 192.205 ;
        RECT 70.320 190.375 70.550 191.365 ;
        RECT 71.245 191.325 71.905 191.525 ;
        RECT 72.075 191.355 74.295 191.525 ;
        RECT 70.720 190.545 71.070 191.195 ;
        RECT 71.245 190.395 71.415 191.325 ;
        RECT 72.075 191.155 72.245 191.355 ;
        RECT 71.585 190.985 72.245 191.155 ;
        RECT 72.415 191.015 73.955 191.185 ;
        RECT 71.585 190.565 71.755 190.985 ;
        RECT 72.415 190.815 72.585 191.015 ;
        RECT 71.985 190.645 72.585 190.815 ;
        RECT 72.755 190.645 73.450 190.845 ;
        RECT 73.710 190.565 73.955 191.015 ;
        RECT 72.075 190.395 72.985 190.475 ;
        RECT 70.320 190.205 71.070 190.375 ;
        RECT 70.315 189.655 70.645 190.035 ;
        RECT 70.815 189.915 71.070 190.205 ;
        RECT 71.245 189.915 71.565 190.395 ;
        RECT 71.735 190.305 72.985 190.395 ;
        RECT 71.735 190.225 72.245 190.305 ;
        RECT 71.735 189.825 71.965 190.225 ;
        RECT 72.135 189.655 72.485 190.045 ;
        RECT 72.655 189.825 72.985 190.305 ;
        RECT 73.155 189.655 73.325 190.475 ;
        RECT 74.125 190.395 74.295 191.355 ;
        RECT 74.465 191.115 75.675 192.205 ;
        RECT 74.465 190.575 74.985 191.115 ;
        RECT 75.845 191.040 76.135 192.205 ;
        RECT 76.305 191.065 76.565 192.205 ;
        RECT 76.735 191.235 77.065 192.035 ;
        RECT 77.235 191.405 77.405 192.205 ;
        RECT 77.605 191.235 77.935 192.035 ;
        RECT 78.135 191.405 78.415 192.205 ;
        RECT 76.735 191.065 78.015 191.235 ;
        RECT 75.155 190.405 75.675 190.945 ;
        RECT 76.330 190.565 76.615 190.895 ;
        RECT 76.815 190.565 77.195 190.895 ;
        RECT 77.365 190.565 77.675 190.895 ;
        RECT 73.830 189.850 74.295 190.395 ;
        RECT 74.465 189.655 75.675 190.405 ;
        RECT 75.845 189.655 76.135 190.380 ;
        RECT 76.310 189.655 76.645 190.395 ;
        RECT 76.815 189.870 77.030 190.565 ;
        RECT 77.365 190.395 77.570 190.565 ;
        RECT 77.845 190.395 78.015 191.065 ;
        RECT 78.195 190.565 78.435 191.235 ;
        RECT 79.525 191.115 83.035 192.205 ;
        RECT 83.580 191.225 83.835 191.895 ;
        RECT 84.015 191.405 84.300 192.205 ;
        RECT 84.480 191.485 84.810 191.995 ;
        RECT 79.525 190.595 81.215 191.115 ;
        RECT 81.385 190.425 83.035 190.945 ;
        RECT 77.220 189.870 77.570 190.395 ;
        RECT 77.740 189.825 78.435 190.395 ;
        RECT 79.525 189.655 83.035 190.425 ;
        RECT 83.580 190.365 83.760 191.225 ;
        RECT 84.480 190.895 84.730 191.485 ;
        RECT 85.080 191.335 85.250 191.945 ;
        RECT 85.420 191.515 85.750 192.205 ;
        RECT 85.980 191.655 86.220 191.945 ;
        RECT 86.420 191.825 86.840 192.205 ;
        RECT 87.020 191.735 87.650 191.985 ;
        RECT 88.120 191.825 88.450 192.205 ;
        RECT 87.020 191.655 87.190 191.735 ;
        RECT 88.620 191.655 88.790 191.945 ;
        RECT 88.970 191.825 89.350 192.205 ;
        RECT 89.590 191.820 90.420 191.990 ;
        RECT 85.980 191.485 87.190 191.655 ;
        RECT 83.930 190.565 84.730 190.895 ;
        RECT 83.580 190.165 83.835 190.365 ;
        RECT 83.495 189.995 83.835 190.165 ;
        RECT 83.580 189.835 83.835 189.995 ;
        RECT 84.015 189.655 84.300 190.115 ;
        RECT 84.480 189.915 84.730 190.565 ;
        RECT 84.930 191.315 85.250 191.335 ;
        RECT 84.930 191.145 86.850 191.315 ;
        RECT 84.930 190.250 85.120 191.145 ;
        RECT 87.020 190.975 87.190 191.485 ;
        RECT 87.360 191.225 87.880 191.535 ;
        RECT 85.290 190.805 87.190 190.975 ;
        RECT 85.290 190.745 85.620 190.805 ;
        RECT 85.770 190.575 86.100 190.635 ;
        RECT 85.440 190.305 86.100 190.575 ;
        RECT 84.930 189.920 85.250 190.250 ;
        RECT 85.430 189.655 86.090 190.135 ;
        RECT 86.290 190.045 86.460 190.805 ;
        RECT 87.360 190.635 87.540 191.045 ;
        RECT 86.630 190.465 86.960 190.585 ;
        RECT 87.710 190.465 87.880 191.225 ;
        RECT 86.630 190.295 87.880 190.465 ;
        RECT 88.050 191.405 89.420 191.655 ;
        RECT 88.050 190.635 88.240 191.405 ;
        RECT 89.170 191.145 89.420 191.405 ;
        RECT 88.410 190.975 88.660 191.135 ;
        RECT 89.590 190.975 89.760 191.820 ;
        RECT 90.655 191.535 90.825 192.035 ;
        RECT 90.995 191.705 91.325 192.205 ;
        RECT 89.930 191.145 90.430 191.525 ;
        RECT 90.655 191.365 91.350 191.535 ;
        RECT 88.410 190.805 89.760 190.975 ;
        RECT 89.340 190.765 89.760 190.805 ;
        RECT 88.050 190.295 88.470 190.635 ;
        RECT 88.760 190.305 89.170 190.635 ;
        RECT 86.290 189.875 87.140 190.045 ;
        RECT 87.700 189.655 88.020 190.115 ;
        RECT 88.220 189.865 88.470 190.295 ;
        RECT 88.760 189.655 89.170 190.095 ;
        RECT 89.340 190.035 89.510 190.765 ;
        RECT 89.680 190.215 90.030 190.585 ;
        RECT 90.210 190.275 90.430 191.145 ;
        RECT 90.600 190.575 91.010 191.195 ;
        RECT 91.180 190.395 91.350 191.365 ;
        RECT 90.655 190.205 91.350 190.395 ;
        RECT 89.340 189.835 90.355 190.035 ;
        RECT 90.655 189.875 90.825 190.205 ;
        RECT 90.995 189.655 91.325 190.035 ;
        RECT 91.540 189.915 91.765 192.035 ;
        RECT 91.935 191.705 92.265 192.205 ;
        RECT 92.435 191.535 92.605 192.035 ;
        RECT 91.940 191.365 92.605 191.535 ;
        RECT 91.940 190.375 92.170 191.365 ;
        RECT 92.955 191.275 93.125 192.035 ;
        RECT 93.305 191.445 93.635 192.205 ;
        RECT 92.340 190.545 92.690 191.195 ;
        RECT 92.955 191.105 93.620 191.275 ;
        RECT 93.805 191.130 94.075 192.035 ;
        RECT 94.245 191.370 94.630 192.205 ;
        RECT 94.800 191.200 95.060 192.005 ;
        RECT 95.230 191.370 95.490 192.205 ;
        RECT 95.660 191.200 95.915 192.005 ;
        RECT 96.090 191.370 96.350 192.205 ;
        RECT 96.520 191.200 96.775 192.005 ;
        RECT 96.950 191.370 97.295 192.205 ;
        RECT 97.465 191.445 97.980 191.855 ;
        RECT 98.215 191.445 98.385 192.205 ;
        RECT 98.555 191.865 100.585 192.035 ;
        RECT 93.450 190.960 93.620 191.105 ;
        RECT 92.885 190.555 93.215 190.925 ;
        RECT 93.450 190.630 93.735 190.960 ;
        RECT 93.450 190.375 93.620 190.630 ;
        RECT 91.940 190.205 92.605 190.375 ;
        RECT 91.935 189.655 92.265 190.035 ;
        RECT 92.435 189.915 92.605 190.205 ;
        RECT 92.955 190.205 93.620 190.375 ;
        RECT 93.905 190.330 94.075 191.130 ;
        RECT 92.955 189.825 93.125 190.205 ;
        RECT 93.305 189.655 93.635 190.035 ;
        RECT 93.815 189.825 94.075 190.330 ;
        RECT 94.245 191.030 97.275 191.200 ;
        RECT 94.245 190.465 94.545 191.030 ;
        RECT 94.720 190.635 96.935 190.860 ;
        RECT 97.105 190.465 97.275 191.030 ;
        RECT 97.465 190.635 97.805 191.445 ;
        RECT 98.555 191.200 98.725 191.865 ;
        RECT 99.120 191.525 100.245 191.695 ;
        RECT 97.975 191.010 98.725 191.200 ;
        RECT 98.895 191.185 99.905 191.355 ;
        RECT 97.465 190.465 98.695 190.635 ;
        RECT 94.245 190.295 97.275 190.465 ;
        RECT 94.765 189.655 95.065 190.125 ;
        RECT 95.235 189.850 95.490 190.295 ;
        RECT 95.660 189.655 95.920 190.125 ;
        RECT 96.090 189.850 96.350 190.295 ;
        RECT 96.520 189.655 96.815 190.125 ;
        RECT 97.740 189.860 97.985 190.465 ;
        RECT 98.205 189.655 98.715 190.190 ;
        RECT 98.895 189.825 99.085 191.185 ;
        RECT 99.255 190.845 99.530 190.985 ;
        RECT 99.255 190.675 99.535 190.845 ;
        RECT 99.255 189.825 99.530 190.675 ;
        RECT 99.735 190.385 99.905 191.185 ;
        RECT 100.075 190.395 100.245 191.525 ;
        RECT 100.415 190.895 100.585 191.865 ;
        RECT 100.755 191.065 100.925 192.205 ;
        RECT 101.095 191.065 101.430 192.035 ;
        RECT 100.415 190.565 100.610 190.895 ;
        RECT 100.835 190.565 101.090 190.895 ;
        RECT 100.835 190.395 101.005 190.565 ;
        RECT 101.260 190.395 101.430 191.065 ;
        RECT 101.605 191.040 101.895 192.205 ;
        RECT 102.155 191.275 102.325 192.035 ;
        RECT 102.505 191.445 102.835 192.205 ;
        RECT 102.155 191.105 102.820 191.275 ;
        RECT 103.005 191.130 103.275 192.035 ;
        RECT 102.650 190.960 102.820 191.105 ;
        RECT 102.085 190.555 102.415 190.925 ;
        RECT 102.650 190.630 102.935 190.960 ;
        RECT 100.075 190.225 101.005 190.395 ;
        RECT 100.075 190.190 100.250 190.225 ;
        RECT 99.720 189.825 100.250 190.190 ;
        RECT 100.675 189.655 101.005 190.055 ;
        RECT 101.175 189.825 101.430 190.395 ;
        RECT 101.605 189.655 101.895 190.380 ;
        RECT 102.650 190.375 102.820 190.630 ;
        RECT 102.155 190.205 102.820 190.375 ;
        RECT 103.105 190.330 103.275 191.130 ;
        RECT 103.445 191.115 104.655 192.205 ;
        RECT 104.825 191.445 105.340 191.855 ;
        RECT 105.575 191.445 105.745 192.205 ;
        RECT 105.915 191.865 107.945 192.035 ;
        RECT 103.445 190.575 103.965 191.115 ;
        RECT 104.135 190.405 104.655 190.945 ;
        RECT 104.825 190.635 105.165 191.445 ;
        RECT 105.915 191.200 106.085 191.865 ;
        RECT 106.480 191.525 107.605 191.695 ;
        RECT 105.335 191.010 106.085 191.200 ;
        RECT 106.255 191.185 107.265 191.355 ;
        RECT 104.825 190.465 106.055 190.635 ;
        RECT 102.155 189.825 102.325 190.205 ;
        RECT 102.505 189.655 102.835 190.035 ;
        RECT 103.015 189.825 103.275 190.330 ;
        RECT 103.445 189.655 104.655 190.405 ;
        RECT 105.100 189.860 105.345 190.465 ;
        RECT 105.565 189.655 106.075 190.190 ;
        RECT 106.255 189.825 106.445 191.185 ;
        RECT 106.615 190.845 106.890 190.985 ;
        RECT 106.615 190.675 106.895 190.845 ;
        RECT 106.615 189.825 106.890 190.675 ;
        RECT 107.095 190.385 107.265 191.185 ;
        RECT 107.435 190.395 107.605 191.525 ;
        RECT 107.775 190.895 107.945 191.865 ;
        RECT 108.115 191.065 108.285 192.205 ;
        RECT 108.455 191.065 108.790 192.035 ;
        RECT 107.775 190.565 107.970 190.895 ;
        RECT 108.195 190.565 108.450 190.895 ;
        RECT 108.195 190.395 108.365 190.565 ;
        RECT 108.620 190.395 108.790 191.065 ;
        RECT 107.435 190.225 108.365 190.395 ;
        RECT 107.435 190.190 107.610 190.225 ;
        RECT 107.080 189.825 107.610 190.190 ;
        RECT 108.035 189.655 108.365 190.055 ;
        RECT 108.535 189.825 108.790 190.395 ;
        RECT 108.970 191.015 109.225 191.895 ;
        RECT 109.395 191.065 109.700 192.205 ;
        RECT 110.040 191.825 110.370 192.205 ;
        RECT 110.550 191.655 110.720 191.945 ;
        RECT 110.890 191.745 111.140 192.205 ;
        RECT 109.920 191.485 110.720 191.655 ;
        RECT 111.310 191.695 112.180 192.035 ;
        RECT 108.970 190.365 109.180 191.015 ;
        RECT 109.920 190.895 110.090 191.485 ;
        RECT 111.310 191.315 111.480 191.695 ;
        RECT 112.415 191.575 112.585 192.035 ;
        RECT 112.755 191.745 113.125 192.205 ;
        RECT 113.420 191.605 113.590 191.945 ;
        RECT 113.760 191.775 114.090 192.205 ;
        RECT 114.325 191.605 114.495 191.945 ;
        RECT 110.260 191.145 111.480 191.315 ;
        RECT 111.650 191.235 112.110 191.525 ;
        RECT 112.415 191.405 112.975 191.575 ;
        RECT 113.420 191.435 114.495 191.605 ;
        RECT 114.665 191.705 115.345 192.035 ;
        RECT 115.560 191.705 115.810 192.035 ;
        RECT 115.980 191.745 116.230 192.205 ;
        RECT 112.805 191.265 112.975 191.405 ;
        RECT 111.650 191.225 112.615 191.235 ;
        RECT 111.310 191.055 111.480 191.145 ;
        RECT 111.940 191.065 112.615 191.225 ;
        RECT 109.350 190.865 110.090 190.895 ;
        RECT 109.350 190.565 110.265 190.865 ;
        RECT 109.940 190.390 110.265 190.565 ;
        RECT 108.970 189.835 109.225 190.365 ;
        RECT 109.395 189.655 109.700 190.115 ;
        RECT 109.945 190.035 110.265 190.390 ;
        RECT 110.435 190.605 110.975 190.975 ;
        RECT 111.310 190.885 111.715 191.055 ;
        RECT 110.435 190.205 110.675 190.605 ;
        RECT 111.155 190.435 111.375 190.715 ;
        RECT 110.845 190.265 111.375 190.435 ;
        RECT 110.845 190.035 111.015 190.265 ;
        RECT 111.545 190.105 111.715 190.885 ;
        RECT 111.885 190.275 112.235 190.895 ;
        RECT 112.405 190.275 112.615 191.065 ;
        RECT 112.805 191.095 114.305 191.265 ;
        RECT 112.805 190.405 112.975 191.095 ;
        RECT 114.665 190.925 114.835 191.705 ;
        RECT 115.640 191.575 115.810 191.705 ;
        RECT 113.145 190.755 114.835 190.925 ;
        RECT 115.005 191.145 115.470 191.535 ;
        RECT 115.640 191.405 116.035 191.575 ;
        RECT 113.145 190.575 113.315 190.755 ;
        RECT 109.945 189.865 111.015 190.035 ;
        RECT 111.185 189.655 111.375 190.095 ;
        RECT 111.545 189.825 112.495 190.105 ;
        RECT 112.805 190.015 113.065 190.405 ;
        RECT 113.485 190.335 114.275 190.585 ;
        RECT 112.715 189.845 113.065 190.015 ;
        RECT 113.275 189.655 113.605 190.115 ;
        RECT 114.480 190.045 114.650 190.755 ;
        RECT 115.005 190.555 115.175 191.145 ;
        RECT 114.820 190.335 115.175 190.555 ;
        RECT 115.345 190.335 115.695 190.955 ;
        RECT 115.865 190.045 116.035 191.405 ;
        RECT 116.400 191.235 116.725 192.020 ;
        RECT 116.205 190.185 116.665 191.235 ;
        RECT 114.480 189.875 115.335 190.045 ;
        RECT 115.540 189.875 116.035 190.045 ;
        RECT 116.205 189.655 116.535 190.015 ;
        RECT 116.895 189.915 117.065 192.035 ;
        RECT 117.235 191.705 117.565 192.205 ;
        RECT 117.735 191.535 117.990 192.035 ;
        RECT 117.240 191.365 117.990 191.535 ;
        RECT 117.240 190.375 117.470 191.365 ;
        RECT 117.640 190.545 117.990 191.195 ;
        RECT 118.165 191.130 118.435 192.035 ;
        RECT 118.605 191.445 118.935 192.205 ;
        RECT 119.115 191.275 119.285 192.035 ;
        RECT 117.240 190.205 117.990 190.375 ;
        RECT 117.235 189.655 117.565 190.035 ;
        RECT 117.735 189.915 117.990 190.205 ;
        RECT 118.165 190.330 118.335 191.130 ;
        RECT 118.620 191.105 119.285 191.275 ;
        RECT 119.545 191.115 120.755 192.205 ;
        RECT 120.930 191.770 126.275 192.205 ;
        RECT 118.620 190.960 118.790 191.105 ;
        RECT 118.505 190.630 118.790 190.960 ;
        RECT 118.620 190.375 118.790 190.630 ;
        RECT 119.025 190.555 119.355 190.925 ;
        RECT 119.545 190.575 120.065 191.115 ;
        RECT 120.235 190.405 120.755 190.945 ;
        RECT 122.520 190.520 122.870 191.770 ;
        RECT 126.445 191.115 127.655 192.205 ;
        RECT 118.165 189.825 118.425 190.330 ;
        RECT 118.620 190.205 119.285 190.375 ;
        RECT 118.605 189.655 118.935 190.035 ;
        RECT 119.115 189.825 119.285 190.205 ;
        RECT 119.545 189.655 120.755 190.405 ;
        RECT 124.350 190.200 124.690 191.030 ;
        RECT 126.445 190.575 126.965 191.115 ;
        RECT 127.135 190.405 127.655 190.945 ;
        RECT 120.930 189.655 126.275 190.200 ;
        RECT 126.445 189.655 127.655 190.405 ;
        RECT 14.580 189.485 127.740 189.655 ;
        RECT 14.665 188.735 15.875 189.485 ;
        RECT 14.665 188.195 15.185 188.735 ;
        RECT 16.505 188.715 18.175 189.485 ;
        RECT 18.350 188.940 23.695 189.485 ;
        RECT 23.870 188.940 29.215 189.485 ;
        RECT 15.355 188.025 15.875 188.565 ;
        RECT 14.665 186.935 15.875 188.025 ;
        RECT 16.505 188.025 17.255 188.545 ;
        RECT 17.425 188.195 18.175 188.715 ;
        RECT 16.505 186.935 18.175 188.025 ;
        RECT 19.940 187.370 20.290 188.620 ;
        RECT 21.770 188.110 22.110 188.940 ;
        RECT 25.460 187.370 25.810 188.620 ;
        RECT 27.290 188.110 27.630 188.940 ;
        RECT 29.445 188.665 29.655 189.485 ;
        RECT 29.825 188.685 30.155 189.315 ;
        RECT 29.825 188.085 30.075 188.685 ;
        RECT 30.325 188.665 30.555 189.485 ;
        RECT 30.765 188.735 31.975 189.485 ;
        RECT 30.245 188.245 30.575 188.495 ;
        RECT 18.350 186.935 23.695 187.370 ;
        RECT 23.870 186.935 29.215 187.370 ;
        RECT 29.445 186.935 29.655 188.075 ;
        RECT 29.825 187.105 30.155 188.085 ;
        RECT 30.325 186.935 30.555 188.075 ;
        RECT 30.765 188.025 31.285 188.565 ;
        RECT 31.455 188.195 31.975 188.735 ;
        RECT 32.145 188.715 35.655 189.485 ;
        RECT 32.145 188.025 33.835 188.545 ;
        RECT 34.005 188.195 35.655 188.715 ;
        RECT 35.865 188.665 36.095 189.485 ;
        RECT 36.265 188.685 36.595 189.315 ;
        RECT 35.845 188.245 36.175 188.495 ;
        RECT 36.345 188.085 36.595 188.685 ;
        RECT 36.765 188.665 36.975 189.485 ;
        RECT 37.205 188.760 37.495 189.485 ;
        RECT 37.670 188.775 37.925 189.305 ;
        RECT 38.095 189.025 38.400 189.485 ;
        RECT 38.645 189.105 39.715 189.275 ;
        RECT 37.670 188.125 37.880 188.775 ;
        RECT 38.645 188.750 38.965 189.105 ;
        RECT 38.640 188.575 38.965 188.750 ;
        RECT 38.050 188.275 38.965 188.575 ;
        RECT 39.135 188.535 39.375 188.935 ;
        RECT 39.545 188.875 39.715 189.105 ;
        RECT 39.885 189.045 40.075 189.485 ;
        RECT 40.245 189.035 41.195 189.315 ;
        RECT 41.415 189.125 41.765 189.295 ;
        RECT 39.545 188.705 40.075 188.875 ;
        RECT 38.050 188.245 38.790 188.275 ;
        RECT 30.765 186.935 31.975 188.025 ;
        RECT 32.145 186.935 35.655 188.025 ;
        RECT 35.865 186.935 36.095 188.075 ;
        RECT 36.265 187.105 36.595 188.085 ;
        RECT 36.765 186.935 36.975 188.075 ;
        RECT 37.205 186.935 37.495 188.100 ;
        RECT 37.670 187.245 37.925 188.125 ;
        RECT 38.095 186.935 38.400 188.075 ;
        RECT 38.620 187.655 38.790 188.245 ;
        RECT 39.135 188.165 39.675 188.535 ;
        RECT 39.855 188.425 40.075 188.705 ;
        RECT 40.245 188.255 40.415 189.035 ;
        RECT 40.010 188.085 40.415 188.255 ;
        RECT 40.585 188.245 40.935 188.865 ;
        RECT 40.010 187.995 40.180 188.085 ;
        RECT 41.105 188.075 41.315 188.865 ;
        RECT 38.960 187.825 40.180 187.995 ;
        RECT 40.640 187.915 41.315 188.075 ;
        RECT 38.620 187.485 39.420 187.655 ;
        RECT 38.740 186.935 39.070 187.315 ;
        RECT 39.250 187.195 39.420 187.485 ;
        RECT 40.010 187.445 40.180 187.825 ;
        RECT 40.350 187.905 41.315 187.915 ;
        RECT 41.505 188.735 41.765 189.125 ;
        RECT 41.975 189.025 42.305 189.485 ;
        RECT 43.180 189.095 44.035 189.265 ;
        RECT 44.240 189.095 44.735 189.265 ;
        RECT 44.905 189.125 45.235 189.485 ;
        RECT 41.505 188.045 41.675 188.735 ;
        RECT 41.845 188.385 42.015 188.565 ;
        RECT 42.185 188.555 42.975 188.805 ;
        RECT 43.180 188.385 43.350 189.095 ;
        RECT 43.520 188.585 43.875 188.805 ;
        RECT 41.845 188.215 43.535 188.385 ;
        RECT 40.350 187.615 40.810 187.905 ;
        RECT 41.505 187.875 43.005 188.045 ;
        RECT 41.505 187.735 41.675 187.875 ;
        RECT 41.115 187.565 41.675 187.735 ;
        RECT 39.590 186.935 39.840 187.395 ;
        RECT 40.010 187.105 40.880 187.445 ;
        RECT 41.115 187.105 41.285 187.565 ;
        RECT 42.120 187.535 43.195 187.705 ;
        RECT 41.455 186.935 41.825 187.395 ;
        RECT 42.120 187.195 42.290 187.535 ;
        RECT 42.460 186.935 42.790 187.365 ;
        RECT 43.025 187.195 43.195 187.535 ;
        RECT 43.365 187.435 43.535 188.215 ;
        RECT 43.705 187.995 43.875 188.585 ;
        RECT 44.045 188.185 44.395 188.805 ;
        RECT 43.705 187.605 44.170 187.995 ;
        RECT 44.565 187.735 44.735 189.095 ;
        RECT 44.905 187.905 45.365 188.955 ;
        RECT 44.340 187.565 44.735 187.735 ;
        RECT 44.340 187.435 44.510 187.565 ;
        RECT 43.365 187.105 44.045 187.435 ;
        RECT 44.260 187.105 44.510 187.435 ;
        RECT 44.680 186.935 44.930 187.395 ;
        RECT 45.100 187.120 45.425 187.905 ;
        RECT 45.595 187.105 45.765 189.225 ;
        RECT 45.935 189.105 46.265 189.485 ;
        RECT 46.435 188.935 46.690 189.225 ;
        RECT 46.955 189.005 47.255 189.485 ;
        RECT 45.940 188.765 46.690 188.935 ;
        RECT 47.425 188.835 47.685 189.290 ;
        RECT 47.855 189.005 48.115 189.485 ;
        RECT 48.295 188.835 48.555 189.290 ;
        RECT 48.725 189.005 48.975 189.485 ;
        RECT 49.155 188.835 49.415 189.290 ;
        RECT 49.585 189.005 49.835 189.485 ;
        RECT 50.015 188.835 50.275 189.290 ;
        RECT 50.445 189.005 50.690 189.485 ;
        RECT 50.860 188.835 51.135 189.290 ;
        RECT 51.305 189.005 51.550 189.485 ;
        RECT 51.720 188.835 51.980 189.290 ;
        RECT 52.150 189.005 52.410 189.485 ;
        RECT 52.580 188.835 52.840 189.290 ;
        RECT 53.010 189.005 53.270 189.485 ;
        RECT 53.440 188.835 53.700 189.290 ;
        RECT 53.870 188.925 54.130 189.485 ;
        RECT 45.940 187.775 46.170 188.765 ;
        RECT 46.955 188.665 53.700 188.835 ;
        RECT 46.340 187.945 46.690 188.595 ;
        RECT 46.955 188.075 48.120 188.665 ;
        RECT 54.300 188.495 54.550 189.305 ;
        RECT 54.730 188.960 54.990 189.485 ;
        RECT 55.160 188.495 55.410 189.305 ;
        RECT 55.590 188.975 55.895 189.485 ;
        RECT 48.290 188.245 55.410 188.495 ;
        RECT 55.580 188.245 55.895 188.805 ;
        RECT 56.340 188.675 56.585 189.280 ;
        RECT 56.805 188.950 57.315 189.485 ;
        RECT 56.065 188.505 57.295 188.675 ;
        RECT 46.955 187.850 53.700 188.075 ;
        RECT 45.940 187.605 46.690 187.775 ;
        RECT 45.935 186.935 46.265 187.435 ;
        RECT 46.435 187.105 46.690 187.605 ;
        RECT 46.955 186.935 47.225 187.680 ;
        RECT 47.395 187.110 47.685 187.850 ;
        RECT 48.295 187.835 53.700 187.850 ;
        RECT 47.855 186.940 48.110 187.665 ;
        RECT 48.295 187.110 48.555 187.835 ;
        RECT 48.725 186.940 48.970 187.665 ;
        RECT 49.155 187.110 49.415 187.835 ;
        RECT 49.585 186.940 49.830 187.665 ;
        RECT 50.015 187.110 50.275 187.835 ;
        RECT 50.445 186.940 50.690 187.665 ;
        RECT 50.860 187.110 51.120 187.835 ;
        RECT 51.290 186.940 51.550 187.665 ;
        RECT 51.720 187.110 51.980 187.835 ;
        RECT 52.150 186.940 52.410 187.665 ;
        RECT 52.580 187.110 52.840 187.835 ;
        RECT 53.010 186.940 53.270 187.665 ;
        RECT 53.440 187.110 53.700 187.835 ;
        RECT 53.870 186.940 54.130 187.735 ;
        RECT 54.300 187.110 54.550 188.245 ;
        RECT 47.855 186.935 54.130 186.940 ;
        RECT 54.730 186.935 54.990 187.745 ;
        RECT 55.165 187.105 55.410 188.245 ;
        RECT 55.590 186.935 55.885 187.745 ;
        RECT 56.065 187.695 56.405 188.505 ;
        RECT 56.575 187.940 57.325 188.130 ;
        RECT 56.065 187.285 56.580 187.695 ;
        RECT 56.815 186.935 56.985 187.695 ;
        RECT 57.155 187.275 57.325 187.940 ;
        RECT 57.495 187.955 57.685 189.315 ;
        RECT 57.855 189.145 58.130 189.315 ;
        RECT 57.855 188.975 58.135 189.145 ;
        RECT 57.855 188.155 58.130 188.975 ;
        RECT 58.320 188.950 58.850 189.315 ;
        RECT 59.275 189.085 59.605 189.485 ;
        RECT 58.675 188.915 58.850 188.950 ;
        RECT 58.335 187.955 58.505 188.755 ;
        RECT 57.495 187.785 58.505 187.955 ;
        RECT 58.675 188.745 59.605 188.915 ;
        RECT 59.775 188.745 60.030 189.315 ;
        RECT 58.675 187.615 58.845 188.745 ;
        RECT 59.435 188.575 59.605 188.745 ;
        RECT 57.720 187.445 58.845 187.615 ;
        RECT 59.015 188.245 59.210 188.575 ;
        RECT 59.435 188.245 59.690 188.575 ;
        RECT 59.015 187.275 59.185 188.245 ;
        RECT 59.860 188.075 60.030 188.745 ;
        RECT 57.155 187.105 59.185 187.275 ;
        RECT 59.355 186.935 59.525 188.075 ;
        RECT 59.695 187.105 60.030 188.075 ;
        RECT 60.205 188.810 60.465 189.315 ;
        RECT 60.645 189.105 60.975 189.485 ;
        RECT 61.155 188.935 61.325 189.315 ;
        RECT 60.205 188.010 60.375 188.810 ;
        RECT 60.660 188.765 61.325 188.935 ;
        RECT 60.660 188.510 60.830 188.765 ;
        RECT 61.585 188.735 62.795 189.485 ;
        RECT 62.965 188.760 63.255 189.485 ;
        RECT 64.000 188.855 64.285 189.315 ;
        RECT 64.455 189.025 64.725 189.485 ;
        RECT 60.545 188.180 60.830 188.510 ;
        RECT 61.065 188.215 61.395 188.585 ;
        RECT 60.660 188.035 60.830 188.180 ;
        RECT 60.205 187.105 60.475 188.010 ;
        RECT 60.660 187.865 61.325 188.035 ;
        RECT 60.645 186.935 60.975 187.695 ;
        RECT 61.155 187.105 61.325 187.865 ;
        RECT 61.585 188.025 62.105 188.565 ;
        RECT 62.275 188.195 62.795 188.735 ;
        RECT 64.000 188.685 64.955 188.855 ;
        RECT 61.585 186.935 62.795 188.025 ;
        RECT 62.965 186.935 63.255 188.100 ;
        RECT 63.885 187.955 64.575 188.515 ;
        RECT 64.745 187.785 64.955 188.685 ;
        RECT 64.000 187.565 64.955 187.785 ;
        RECT 65.125 188.515 65.525 189.315 ;
        RECT 65.715 188.855 65.995 189.315 ;
        RECT 66.515 189.025 66.840 189.485 ;
        RECT 65.715 188.685 66.840 188.855 ;
        RECT 67.010 188.745 67.395 189.315 ;
        RECT 66.390 188.575 66.840 188.685 ;
        RECT 65.125 187.955 66.220 188.515 ;
        RECT 66.390 188.245 66.945 188.575 ;
        RECT 64.000 187.105 64.285 187.565 ;
        RECT 64.455 186.935 64.725 187.395 ;
        RECT 65.125 187.105 65.525 187.955 ;
        RECT 66.390 187.785 66.840 188.245 ;
        RECT 67.115 188.075 67.395 188.745 ;
        RECT 67.565 188.715 70.155 189.485 ;
        RECT 70.330 188.940 75.675 189.485 ;
        RECT 75.850 188.940 81.195 189.485 ;
        RECT 81.370 188.940 86.715 189.485 ;
        RECT 65.715 187.565 66.840 187.785 ;
        RECT 65.715 187.105 65.995 187.565 ;
        RECT 66.515 186.935 66.840 187.395 ;
        RECT 67.010 187.105 67.395 188.075 ;
        RECT 67.565 188.025 68.775 188.545 ;
        RECT 68.945 188.195 70.155 188.715 ;
        RECT 67.565 186.935 70.155 188.025 ;
        RECT 71.920 187.370 72.270 188.620 ;
        RECT 73.750 188.110 74.090 188.940 ;
        RECT 77.440 187.370 77.790 188.620 ;
        RECT 79.270 188.110 79.610 188.940 ;
        RECT 82.960 187.370 83.310 188.620 ;
        RECT 84.790 188.110 85.130 188.940 ;
        RECT 86.945 188.665 87.155 189.485 ;
        RECT 87.325 188.685 87.655 189.315 ;
        RECT 87.325 188.085 87.575 188.685 ;
        RECT 87.825 188.665 88.055 189.485 ;
        RECT 88.725 188.760 89.015 189.485 ;
        RECT 89.275 188.935 89.445 189.315 ;
        RECT 89.625 189.105 89.955 189.485 ;
        RECT 89.275 188.765 89.940 188.935 ;
        RECT 90.135 188.810 90.395 189.315 ;
        RECT 87.745 188.245 88.075 188.495 ;
        RECT 89.205 188.215 89.535 188.585 ;
        RECT 89.770 188.510 89.940 188.765 ;
        RECT 89.770 188.180 90.055 188.510 ;
        RECT 70.330 186.935 75.675 187.370 ;
        RECT 75.850 186.935 81.195 187.370 ;
        RECT 81.370 186.935 86.715 187.370 ;
        RECT 86.945 186.935 87.155 188.075 ;
        RECT 87.325 187.105 87.655 188.085 ;
        RECT 87.825 186.935 88.055 188.075 ;
        RECT 88.725 186.935 89.015 188.100 ;
        RECT 89.770 188.035 89.940 188.180 ;
        RECT 89.275 187.865 89.940 188.035 ;
        RECT 90.225 188.010 90.395 188.810 ;
        RECT 90.565 188.715 92.235 189.485 ;
        RECT 92.410 188.940 97.755 189.485 ;
        RECT 89.275 187.105 89.445 187.865 ;
        RECT 89.625 186.935 89.955 187.695 ;
        RECT 90.125 187.105 90.395 188.010 ;
        RECT 90.565 188.025 91.315 188.545 ;
        RECT 91.485 188.195 92.235 188.715 ;
        RECT 90.565 186.935 92.235 188.025 ;
        RECT 94.000 187.370 94.350 188.620 ;
        RECT 95.830 188.110 96.170 188.940 ;
        RECT 97.930 188.775 98.185 189.305 ;
        RECT 98.355 189.025 98.660 189.485 ;
        RECT 98.905 189.105 99.975 189.275 ;
        RECT 97.930 188.125 98.140 188.775 ;
        RECT 98.905 188.750 99.225 189.105 ;
        RECT 98.900 188.575 99.225 188.750 ;
        RECT 98.310 188.275 99.225 188.575 ;
        RECT 99.395 188.535 99.635 188.935 ;
        RECT 99.805 188.875 99.975 189.105 ;
        RECT 100.145 189.045 100.335 189.485 ;
        RECT 100.505 189.035 101.455 189.315 ;
        RECT 101.675 189.125 102.025 189.295 ;
        RECT 99.805 188.705 100.335 188.875 ;
        RECT 98.310 188.245 99.050 188.275 ;
        RECT 92.410 186.935 97.755 187.370 ;
        RECT 97.930 187.245 98.185 188.125 ;
        RECT 98.355 186.935 98.660 188.075 ;
        RECT 98.880 187.655 99.050 188.245 ;
        RECT 99.395 188.165 99.935 188.535 ;
        RECT 100.115 188.425 100.335 188.705 ;
        RECT 100.505 188.255 100.675 189.035 ;
        RECT 100.270 188.085 100.675 188.255 ;
        RECT 100.845 188.245 101.195 188.865 ;
        RECT 100.270 187.995 100.440 188.085 ;
        RECT 101.365 188.075 101.575 188.865 ;
        RECT 99.220 187.825 100.440 187.995 ;
        RECT 100.900 187.915 101.575 188.075 ;
        RECT 98.880 187.485 99.680 187.655 ;
        RECT 99.000 186.935 99.330 187.315 ;
        RECT 99.510 187.195 99.680 187.485 ;
        RECT 100.270 187.445 100.440 187.825 ;
        RECT 100.610 187.905 101.575 187.915 ;
        RECT 101.765 188.735 102.025 189.125 ;
        RECT 102.235 189.025 102.565 189.485 ;
        RECT 103.440 189.095 104.295 189.265 ;
        RECT 104.500 189.095 104.995 189.265 ;
        RECT 105.165 189.125 105.495 189.485 ;
        RECT 101.765 188.045 101.935 188.735 ;
        RECT 102.105 188.385 102.275 188.565 ;
        RECT 102.445 188.555 103.235 188.805 ;
        RECT 103.440 188.385 103.610 189.095 ;
        RECT 103.780 188.585 104.135 188.805 ;
        RECT 102.105 188.215 103.795 188.385 ;
        RECT 100.610 187.615 101.070 187.905 ;
        RECT 101.765 187.875 103.265 188.045 ;
        RECT 101.765 187.735 101.935 187.875 ;
        RECT 101.375 187.565 101.935 187.735 ;
        RECT 99.850 186.935 100.100 187.395 ;
        RECT 100.270 187.105 101.140 187.445 ;
        RECT 101.375 187.105 101.545 187.565 ;
        RECT 102.380 187.535 103.455 187.705 ;
        RECT 101.715 186.935 102.085 187.395 ;
        RECT 102.380 187.195 102.550 187.535 ;
        RECT 102.720 186.935 103.050 187.365 ;
        RECT 103.285 187.195 103.455 187.535 ;
        RECT 103.625 187.435 103.795 188.215 ;
        RECT 103.965 187.995 104.135 188.585 ;
        RECT 104.305 188.185 104.655 188.805 ;
        RECT 103.965 187.605 104.430 187.995 ;
        RECT 104.825 187.735 104.995 189.095 ;
        RECT 105.165 187.905 105.625 188.955 ;
        RECT 104.600 187.565 104.995 187.735 ;
        RECT 104.600 187.435 104.770 187.565 ;
        RECT 103.625 187.105 104.305 187.435 ;
        RECT 104.520 187.105 104.770 187.435 ;
        RECT 104.940 186.935 105.190 187.395 ;
        RECT 105.360 187.120 105.685 187.905 ;
        RECT 105.855 187.105 106.025 189.225 ;
        RECT 106.195 189.105 106.525 189.485 ;
        RECT 106.695 188.935 106.950 189.225 ;
        RECT 106.200 188.765 106.950 188.935 ;
        RECT 106.200 187.775 106.430 188.765 ;
        RECT 107.125 188.745 107.510 189.315 ;
        RECT 107.680 189.025 108.005 189.485 ;
        RECT 108.525 188.855 108.805 189.315 ;
        RECT 106.600 187.945 106.950 188.595 ;
        RECT 107.125 188.075 107.405 188.745 ;
        RECT 107.680 188.685 108.805 188.855 ;
        RECT 107.680 188.575 108.130 188.685 ;
        RECT 107.575 188.245 108.130 188.575 ;
        RECT 108.995 188.515 109.395 189.315 ;
        RECT 109.795 189.025 110.065 189.485 ;
        RECT 110.235 188.855 110.520 189.315 ;
        RECT 106.200 187.605 106.950 187.775 ;
        RECT 106.195 186.935 106.525 187.435 ;
        RECT 106.695 187.105 106.950 187.605 ;
        RECT 107.125 187.105 107.510 188.075 ;
        RECT 107.680 187.785 108.130 188.245 ;
        RECT 108.300 187.955 109.395 188.515 ;
        RECT 107.680 187.565 108.805 187.785 ;
        RECT 107.680 186.935 108.005 187.395 ;
        RECT 108.525 187.105 108.805 187.565 ;
        RECT 108.995 187.105 109.395 187.955 ;
        RECT 109.565 188.685 110.520 188.855 ;
        RECT 111.265 188.715 112.935 189.485 ;
        RECT 113.195 188.935 113.365 189.315 ;
        RECT 113.545 189.105 113.875 189.485 ;
        RECT 113.195 188.765 113.860 188.935 ;
        RECT 114.055 188.810 114.315 189.315 ;
        RECT 109.565 187.785 109.775 188.685 ;
        RECT 109.945 187.955 110.635 188.515 ;
        RECT 111.265 188.025 112.015 188.545 ;
        RECT 112.185 188.195 112.935 188.715 ;
        RECT 113.125 188.215 113.455 188.585 ;
        RECT 113.690 188.510 113.860 188.765 ;
        RECT 113.690 188.180 113.975 188.510 ;
        RECT 113.690 188.035 113.860 188.180 ;
        RECT 109.565 187.565 110.520 187.785 ;
        RECT 109.795 186.935 110.065 187.395 ;
        RECT 110.235 187.105 110.520 187.565 ;
        RECT 111.265 186.935 112.935 188.025 ;
        RECT 113.195 187.865 113.860 188.035 ;
        RECT 114.145 188.010 114.315 188.810 ;
        RECT 114.485 188.760 114.775 189.485 ;
        RECT 115.410 188.940 120.755 189.485 ;
        RECT 120.930 188.940 126.275 189.485 ;
        RECT 113.195 187.105 113.365 187.865 ;
        RECT 113.545 186.935 113.875 187.695 ;
        RECT 114.045 187.105 114.315 188.010 ;
        RECT 114.485 186.935 114.775 188.100 ;
        RECT 117.000 187.370 117.350 188.620 ;
        RECT 118.830 188.110 119.170 188.940 ;
        RECT 122.520 187.370 122.870 188.620 ;
        RECT 124.350 188.110 124.690 188.940 ;
        RECT 126.445 188.735 127.655 189.485 ;
        RECT 126.445 188.025 126.965 188.565 ;
        RECT 127.135 188.195 127.655 188.735 ;
        RECT 115.410 186.935 120.755 187.370 ;
        RECT 120.930 186.935 126.275 187.370 ;
        RECT 126.445 186.935 127.655 188.025 ;
        RECT 14.580 186.765 127.740 186.935 ;
        RECT 14.665 185.675 15.875 186.765 ;
        RECT 14.665 184.965 15.185 185.505 ;
        RECT 15.355 185.135 15.875 185.675 ;
        RECT 16.045 185.675 18.635 186.765 ;
        RECT 18.810 186.330 24.155 186.765 ;
        RECT 16.045 185.155 17.255 185.675 ;
        RECT 17.425 184.985 18.635 185.505 ;
        RECT 20.400 185.080 20.750 186.330 ;
        RECT 24.325 185.600 24.615 186.765 ;
        RECT 24.785 185.675 25.995 186.765 ;
        RECT 14.665 184.215 15.875 184.965 ;
        RECT 16.045 184.215 18.635 184.985 ;
        RECT 22.230 184.760 22.570 185.590 ;
        RECT 24.785 185.135 25.305 185.675 ;
        RECT 26.170 185.575 26.425 186.455 ;
        RECT 26.595 185.625 26.900 186.765 ;
        RECT 27.240 186.385 27.570 186.765 ;
        RECT 27.750 186.215 27.920 186.505 ;
        RECT 28.090 186.305 28.340 186.765 ;
        RECT 27.120 186.045 27.920 186.215 ;
        RECT 28.510 186.255 29.380 186.595 ;
        RECT 25.475 184.965 25.995 185.505 ;
        RECT 18.810 184.215 24.155 184.760 ;
        RECT 24.325 184.215 24.615 184.940 ;
        RECT 24.785 184.215 25.995 184.965 ;
        RECT 26.170 184.925 26.380 185.575 ;
        RECT 27.120 185.455 27.290 186.045 ;
        RECT 28.510 185.875 28.680 186.255 ;
        RECT 29.615 186.135 29.785 186.595 ;
        RECT 29.955 186.305 30.325 186.765 ;
        RECT 30.620 186.165 30.790 186.505 ;
        RECT 30.960 186.335 31.290 186.765 ;
        RECT 31.525 186.165 31.695 186.505 ;
        RECT 27.460 185.705 28.680 185.875 ;
        RECT 28.850 185.795 29.310 186.085 ;
        RECT 29.615 185.965 30.175 186.135 ;
        RECT 30.620 185.995 31.695 186.165 ;
        RECT 31.865 186.265 32.545 186.595 ;
        RECT 32.760 186.265 33.010 186.595 ;
        RECT 33.180 186.305 33.430 186.765 ;
        RECT 30.005 185.825 30.175 185.965 ;
        RECT 28.850 185.785 29.815 185.795 ;
        RECT 28.510 185.615 28.680 185.705 ;
        RECT 29.140 185.625 29.815 185.785 ;
        RECT 26.550 185.425 27.290 185.455 ;
        RECT 26.550 185.125 27.465 185.425 ;
        RECT 27.140 184.950 27.465 185.125 ;
        RECT 26.170 184.395 26.425 184.925 ;
        RECT 26.595 184.215 26.900 184.675 ;
        RECT 27.145 184.595 27.465 184.950 ;
        RECT 27.635 185.165 28.175 185.535 ;
        RECT 28.510 185.445 28.915 185.615 ;
        RECT 27.635 184.765 27.875 185.165 ;
        RECT 28.355 184.995 28.575 185.275 ;
        RECT 28.045 184.825 28.575 184.995 ;
        RECT 28.045 184.595 28.215 184.825 ;
        RECT 28.745 184.665 28.915 185.445 ;
        RECT 29.085 184.835 29.435 185.455 ;
        RECT 29.605 184.835 29.815 185.625 ;
        RECT 30.005 185.655 31.505 185.825 ;
        RECT 30.005 184.965 30.175 185.655 ;
        RECT 31.865 185.485 32.035 186.265 ;
        RECT 32.840 186.135 33.010 186.265 ;
        RECT 30.345 185.315 32.035 185.485 ;
        RECT 32.205 185.705 32.670 186.095 ;
        RECT 32.840 185.965 33.235 186.135 ;
        RECT 30.345 185.135 30.515 185.315 ;
        RECT 27.145 184.425 28.215 184.595 ;
        RECT 28.385 184.215 28.575 184.655 ;
        RECT 28.745 184.385 29.695 184.665 ;
        RECT 30.005 184.575 30.265 184.965 ;
        RECT 30.685 184.895 31.475 185.145 ;
        RECT 29.915 184.405 30.265 184.575 ;
        RECT 30.475 184.215 30.805 184.675 ;
        RECT 31.680 184.605 31.850 185.315 ;
        RECT 32.205 185.115 32.375 185.705 ;
        RECT 32.020 184.895 32.375 185.115 ;
        RECT 32.545 184.895 32.895 185.515 ;
        RECT 33.065 184.605 33.235 185.965 ;
        RECT 33.600 185.795 33.925 186.580 ;
        RECT 33.405 184.745 33.865 185.795 ;
        RECT 31.680 184.435 32.535 184.605 ;
        RECT 32.740 184.435 33.235 184.605 ;
        RECT 33.405 184.215 33.735 184.575 ;
        RECT 34.095 184.475 34.265 186.595 ;
        RECT 34.435 186.265 34.765 186.765 ;
        RECT 34.935 186.095 35.190 186.595 ;
        RECT 34.440 185.925 35.190 186.095 ;
        RECT 34.440 184.935 34.670 185.925 ;
        RECT 34.840 185.105 35.190 185.755 ;
        RECT 35.825 185.675 38.415 186.765 ;
        RECT 35.825 185.155 37.035 185.675 ;
        RECT 38.625 185.625 38.855 186.765 ;
        RECT 39.025 185.615 39.355 186.595 ;
        RECT 39.525 185.625 39.735 186.765 ;
        RECT 39.965 186.005 40.480 186.415 ;
        RECT 40.715 186.005 40.885 186.765 ;
        RECT 41.055 186.425 43.085 186.595 ;
        RECT 37.205 184.985 38.415 185.505 ;
        RECT 38.605 185.205 38.935 185.455 ;
        RECT 34.440 184.765 35.190 184.935 ;
        RECT 34.435 184.215 34.765 184.595 ;
        RECT 34.935 184.475 35.190 184.765 ;
        RECT 35.825 184.215 38.415 184.985 ;
        RECT 38.625 184.215 38.855 185.035 ;
        RECT 39.105 185.015 39.355 185.615 ;
        RECT 39.965 185.195 40.305 186.005 ;
        RECT 41.055 185.760 41.225 186.425 ;
        RECT 41.620 186.085 42.745 186.255 ;
        RECT 40.475 185.570 41.225 185.760 ;
        RECT 41.395 185.745 42.405 185.915 ;
        RECT 39.025 184.385 39.355 185.015 ;
        RECT 39.525 184.215 39.735 185.035 ;
        RECT 39.965 185.025 41.195 185.195 ;
        RECT 40.240 184.420 40.485 185.025 ;
        RECT 40.705 184.215 41.215 184.750 ;
        RECT 41.395 184.385 41.585 185.745 ;
        RECT 41.755 184.725 42.030 185.545 ;
        RECT 42.235 184.945 42.405 185.745 ;
        RECT 42.575 184.955 42.745 186.085 ;
        RECT 42.915 185.455 43.085 186.425 ;
        RECT 43.255 185.625 43.425 186.765 ;
        RECT 43.595 185.625 43.930 186.595 ;
        RECT 42.915 185.125 43.110 185.455 ;
        RECT 43.335 185.125 43.590 185.455 ;
        RECT 43.335 184.955 43.505 185.125 ;
        RECT 43.760 184.955 43.930 185.625 ;
        RECT 42.575 184.785 43.505 184.955 ;
        RECT 42.575 184.750 42.750 184.785 ;
        RECT 41.755 184.555 42.035 184.725 ;
        RECT 41.755 184.385 42.030 184.555 ;
        RECT 42.220 184.385 42.750 184.750 ;
        RECT 43.175 184.215 43.505 184.615 ;
        RECT 43.675 184.385 43.930 184.955 ;
        RECT 44.110 185.625 44.445 186.595 ;
        RECT 44.615 185.625 44.785 186.765 ;
        RECT 44.955 186.425 46.985 186.595 ;
        RECT 44.110 184.955 44.280 185.625 ;
        RECT 44.955 185.455 45.125 186.425 ;
        RECT 44.450 185.125 44.705 185.455 ;
        RECT 44.930 185.125 45.125 185.455 ;
        RECT 45.295 186.085 46.420 186.255 ;
        RECT 44.535 184.955 44.705 185.125 ;
        RECT 45.295 184.955 45.465 186.085 ;
        RECT 44.110 184.385 44.365 184.955 ;
        RECT 44.535 184.785 45.465 184.955 ;
        RECT 45.635 185.745 46.645 185.915 ;
        RECT 45.635 184.945 45.805 185.745 ;
        RECT 45.290 184.750 45.465 184.785 ;
        RECT 44.535 184.215 44.865 184.615 ;
        RECT 45.290 184.385 45.820 184.750 ;
        RECT 46.010 184.725 46.285 185.545 ;
        RECT 46.005 184.555 46.285 184.725 ;
        RECT 46.010 184.385 46.285 184.555 ;
        RECT 46.455 184.385 46.645 185.745 ;
        RECT 46.815 185.760 46.985 186.425 ;
        RECT 47.155 186.005 47.325 186.765 ;
        RECT 47.560 186.005 48.075 186.415 ;
        RECT 46.815 185.570 47.565 185.760 ;
        RECT 47.735 185.195 48.075 186.005 ;
        RECT 48.745 185.625 48.975 186.765 ;
        RECT 49.145 185.615 49.475 186.595 ;
        RECT 49.645 185.625 49.855 186.765 ;
        RECT 48.725 185.205 49.055 185.455 ;
        RECT 46.845 185.025 48.075 185.195 ;
        RECT 46.825 184.215 47.335 184.750 ;
        RECT 47.555 184.420 47.800 185.025 ;
        RECT 48.745 184.215 48.975 185.035 ;
        RECT 49.225 185.015 49.475 185.615 ;
        RECT 50.085 185.600 50.375 186.765 ;
        RECT 50.550 185.575 50.805 186.455 ;
        RECT 50.975 185.625 51.280 186.765 ;
        RECT 51.620 186.385 51.950 186.765 ;
        RECT 52.130 186.215 52.300 186.505 ;
        RECT 52.470 186.305 52.720 186.765 ;
        RECT 51.500 186.045 52.300 186.215 ;
        RECT 52.890 186.255 53.760 186.595 ;
        RECT 49.145 184.385 49.475 185.015 ;
        RECT 49.645 184.215 49.855 185.035 ;
        RECT 50.085 184.215 50.375 184.940 ;
        RECT 50.550 184.925 50.760 185.575 ;
        RECT 51.500 185.455 51.670 186.045 ;
        RECT 52.890 185.875 53.060 186.255 ;
        RECT 53.995 186.135 54.165 186.595 ;
        RECT 54.335 186.305 54.705 186.765 ;
        RECT 55.000 186.165 55.170 186.505 ;
        RECT 55.340 186.335 55.670 186.765 ;
        RECT 55.905 186.165 56.075 186.505 ;
        RECT 51.840 185.705 53.060 185.875 ;
        RECT 53.230 185.795 53.690 186.085 ;
        RECT 53.995 185.965 54.555 186.135 ;
        RECT 55.000 185.995 56.075 186.165 ;
        RECT 56.245 186.265 56.925 186.595 ;
        RECT 57.140 186.265 57.390 186.595 ;
        RECT 57.560 186.305 57.810 186.765 ;
        RECT 54.385 185.825 54.555 185.965 ;
        RECT 53.230 185.785 54.195 185.795 ;
        RECT 52.890 185.615 53.060 185.705 ;
        RECT 53.520 185.625 54.195 185.785 ;
        RECT 50.930 185.425 51.670 185.455 ;
        RECT 50.930 185.125 51.845 185.425 ;
        RECT 51.520 184.950 51.845 185.125 ;
        RECT 50.550 184.395 50.805 184.925 ;
        RECT 50.975 184.215 51.280 184.675 ;
        RECT 51.525 184.595 51.845 184.950 ;
        RECT 52.015 185.165 52.555 185.535 ;
        RECT 52.890 185.445 53.295 185.615 ;
        RECT 52.015 184.765 52.255 185.165 ;
        RECT 52.735 184.995 52.955 185.275 ;
        RECT 52.425 184.825 52.955 184.995 ;
        RECT 52.425 184.595 52.595 184.825 ;
        RECT 53.125 184.665 53.295 185.445 ;
        RECT 53.465 184.835 53.815 185.455 ;
        RECT 53.985 184.835 54.195 185.625 ;
        RECT 54.385 185.655 55.885 185.825 ;
        RECT 54.385 184.965 54.555 185.655 ;
        RECT 56.245 185.485 56.415 186.265 ;
        RECT 57.220 186.135 57.390 186.265 ;
        RECT 54.725 185.315 56.415 185.485 ;
        RECT 56.585 185.705 57.050 186.095 ;
        RECT 57.220 185.965 57.615 186.135 ;
        RECT 54.725 185.135 54.895 185.315 ;
        RECT 51.525 184.425 52.595 184.595 ;
        RECT 52.765 184.215 52.955 184.655 ;
        RECT 53.125 184.385 54.075 184.665 ;
        RECT 54.385 184.575 54.645 184.965 ;
        RECT 55.065 184.895 55.855 185.145 ;
        RECT 54.295 184.405 54.645 184.575 ;
        RECT 54.855 184.215 55.185 184.675 ;
        RECT 56.060 184.605 56.230 185.315 ;
        RECT 56.585 185.115 56.755 185.705 ;
        RECT 56.400 184.895 56.755 185.115 ;
        RECT 56.925 184.895 57.275 185.515 ;
        RECT 57.445 184.605 57.615 185.965 ;
        RECT 57.980 185.795 58.305 186.580 ;
        RECT 57.785 184.745 58.245 185.795 ;
        RECT 56.060 184.435 56.915 184.605 ;
        RECT 57.120 184.435 57.615 184.605 ;
        RECT 57.785 184.215 58.115 184.575 ;
        RECT 58.475 184.475 58.645 186.595 ;
        RECT 58.815 186.265 59.145 186.765 ;
        RECT 59.315 186.095 59.570 186.595 ;
        RECT 60.210 186.330 65.555 186.765 ;
        RECT 65.730 186.330 71.075 186.765 ;
        RECT 58.820 185.925 59.570 186.095 ;
        RECT 58.820 184.935 59.050 185.925 ;
        RECT 59.220 185.105 59.570 185.755 ;
        RECT 61.800 185.080 62.150 186.330 ;
        RECT 58.820 184.765 59.570 184.935 ;
        RECT 58.815 184.215 59.145 184.595 ;
        RECT 59.315 184.475 59.570 184.765 ;
        RECT 63.630 184.760 63.970 185.590 ;
        RECT 67.320 185.080 67.670 186.330 ;
        RECT 69.150 184.760 69.490 185.590 ;
        RECT 60.210 184.215 65.555 184.760 ;
        RECT 65.730 184.215 71.075 184.760 ;
        RECT 71.245 184.385 71.505 186.595 ;
        RECT 71.675 186.385 72.005 186.765 ;
        RECT 72.430 186.215 72.600 186.595 ;
        RECT 72.860 186.385 73.190 186.765 ;
        RECT 73.385 186.215 73.555 186.595 ;
        RECT 73.765 186.385 74.095 186.765 ;
        RECT 74.345 186.215 74.535 186.595 ;
        RECT 74.775 186.385 75.105 186.765 ;
        RECT 75.415 186.265 75.675 186.595 ;
        RECT 71.675 186.045 73.625 186.215 ;
        RECT 71.675 185.125 71.845 186.045 ;
        RECT 72.215 185.455 72.410 185.765 ;
        RECT 72.680 185.455 72.865 185.765 ;
        RECT 72.155 185.125 72.410 185.455 ;
        RECT 72.635 185.125 72.865 185.455 ;
        RECT 71.675 184.215 72.005 184.595 ;
        RECT 72.215 184.550 72.410 185.125 ;
        RECT 72.680 184.545 72.865 185.125 ;
        RECT 73.115 184.555 73.285 185.455 ;
        RECT 73.455 185.055 73.625 186.045 ;
        RECT 73.795 186.045 74.535 186.215 ;
        RECT 73.795 185.535 73.965 186.045 ;
        RECT 74.135 185.705 74.715 185.875 ;
        RECT 74.985 185.755 75.335 186.085 ;
        RECT 74.545 185.585 74.715 185.705 ;
        RECT 75.505 185.585 75.675 186.265 ;
        RECT 75.845 185.600 76.135 186.765 ;
        RECT 76.305 185.675 78.895 186.765 ;
        RECT 79.070 186.330 84.415 186.765 ;
        RECT 73.795 185.365 74.365 185.535 ;
        RECT 74.545 185.415 75.675 185.585 ;
        RECT 73.455 184.725 74.005 185.055 ;
        RECT 74.195 184.885 74.365 185.365 ;
        RECT 74.535 185.075 75.155 185.245 ;
        RECT 74.945 184.895 75.155 185.075 ;
        RECT 74.195 184.555 74.595 184.885 ;
        RECT 75.505 184.715 75.675 185.415 ;
        RECT 76.305 185.155 77.515 185.675 ;
        RECT 77.685 184.985 78.895 185.505 ;
        RECT 80.660 185.080 81.010 186.330 ;
        RECT 84.585 186.005 85.100 186.415 ;
        RECT 85.335 186.005 85.505 186.765 ;
        RECT 85.675 186.425 87.705 186.595 ;
        RECT 73.115 184.385 74.595 184.555 ;
        RECT 74.775 184.215 75.105 184.595 ;
        RECT 75.415 184.385 75.675 184.715 ;
        RECT 75.845 184.215 76.135 184.940 ;
        RECT 76.305 184.215 78.895 184.985 ;
        RECT 82.490 184.760 82.830 185.590 ;
        RECT 84.585 185.195 84.925 186.005 ;
        RECT 85.675 185.760 85.845 186.425 ;
        RECT 86.240 186.085 87.365 186.255 ;
        RECT 85.095 185.570 85.845 185.760 ;
        RECT 86.015 185.745 87.025 185.915 ;
        RECT 84.585 185.025 85.815 185.195 ;
        RECT 79.070 184.215 84.415 184.760 ;
        RECT 84.860 184.420 85.105 185.025 ;
        RECT 85.325 184.215 85.835 184.750 ;
        RECT 86.015 184.385 86.205 185.745 ;
        RECT 86.375 184.725 86.650 185.545 ;
        RECT 86.855 184.945 87.025 185.745 ;
        RECT 87.195 184.955 87.365 186.085 ;
        RECT 87.535 185.455 87.705 186.425 ;
        RECT 87.875 185.625 88.045 186.765 ;
        RECT 88.215 185.625 88.550 186.595 ;
        RECT 88.730 186.330 94.075 186.765 ;
        RECT 87.535 185.125 87.730 185.455 ;
        RECT 87.955 185.125 88.210 185.455 ;
        RECT 87.955 184.955 88.125 185.125 ;
        RECT 88.380 184.955 88.550 185.625 ;
        RECT 90.320 185.080 90.670 186.330 ;
        RECT 94.360 186.135 94.645 186.595 ;
        RECT 94.815 186.305 95.085 186.765 ;
        RECT 94.360 185.915 95.315 186.135 ;
        RECT 87.195 184.785 88.125 184.955 ;
        RECT 87.195 184.750 87.370 184.785 ;
        RECT 86.375 184.555 86.655 184.725 ;
        RECT 86.375 184.385 86.650 184.555 ;
        RECT 86.840 184.385 87.370 184.750 ;
        RECT 87.795 184.215 88.125 184.615 ;
        RECT 88.295 184.385 88.550 184.955 ;
        RECT 92.150 184.760 92.490 185.590 ;
        RECT 94.245 185.185 94.935 185.745 ;
        RECT 95.105 185.015 95.315 185.915 ;
        RECT 94.360 184.845 95.315 185.015 ;
        RECT 95.485 185.745 95.885 186.595 ;
        RECT 96.075 186.135 96.355 186.595 ;
        RECT 96.875 186.305 97.200 186.765 ;
        RECT 96.075 185.915 97.200 186.135 ;
        RECT 95.485 185.185 96.580 185.745 ;
        RECT 96.750 185.455 97.200 185.915 ;
        RECT 97.370 185.625 97.755 186.595 ;
        RECT 98.935 185.835 99.105 186.595 ;
        RECT 99.285 186.005 99.615 186.765 ;
        RECT 98.935 185.665 99.600 185.835 ;
        RECT 99.785 185.690 100.055 186.595 ;
        RECT 88.730 184.215 94.075 184.760 ;
        RECT 94.360 184.385 94.645 184.845 ;
        RECT 94.815 184.215 95.085 184.675 ;
        RECT 95.485 184.385 95.885 185.185 ;
        RECT 96.750 185.125 97.305 185.455 ;
        RECT 96.750 185.015 97.200 185.125 ;
        RECT 96.075 184.845 97.200 185.015 ;
        RECT 97.475 184.955 97.755 185.625 ;
        RECT 99.430 185.520 99.600 185.665 ;
        RECT 98.865 185.115 99.195 185.485 ;
        RECT 99.430 185.190 99.715 185.520 ;
        RECT 96.075 184.385 96.355 184.845 ;
        RECT 96.875 184.215 97.200 184.675 ;
        RECT 97.370 184.385 97.755 184.955 ;
        RECT 99.430 184.935 99.600 185.190 ;
        RECT 98.935 184.765 99.600 184.935 ;
        RECT 99.885 184.890 100.055 185.690 ;
        RECT 100.265 185.625 100.495 186.765 ;
        RECT 100.665 185.615 100.995 186.595 ;
        RECT 101.165 185.625 101.375 186.765 ;
        RECT 100.245 185.205 100.575 185.455 ;
        RECT 98.935 184.385 99.105 184.765 ;
        RECT 99.285 184.215 99.615 184.595 ;
        RECT 99.795 184.385 100.055 184.890 ;
        RECT 100.265 184.215 100.495 185.035 ;
        RECT 100.745 185.015 100.995 185.615 ;
        RECT 101.605 185.600 101.895 186.765 ;
        RECT 102.525 185.625 102.910 186.595 ;
        RECT 103.080 186.305 103.405 186.765 ;
        RECT 103.925 186.135 104.205 186.595 ;
        RECT 103.080 185.915 104.205 186.135 ;
        RECT 100.665 184.385 100.995 185.015 ;
        RECT 101.165 184.215 101.375 185.035 ;
        RECT 102.525 184.955 102.805 185.625 ;
        RECT 103.080 185.455 103.530 185.915 ;
        RECT 104.395 185.745 104.795 186.595 ;
        RECT 105.195 186.305 105.465 186.765 ;
        RECT 105.635 186.135 105.920 186.595 ;
        RECT 102.975 185.125 103.530 185.455 ;
        RECT 103.700 185.185 104.795 185.745 ;
        RECT 103.080 185.015 103.530 185.125 ;
        RECT 101.605 184.215 101.895 184.940 ;
        RECT 102.525 184.385 102.910 184.955 ;
        RECT 103.080 184.845 104.205 185.015 ;
        RECT 103.080 184.215 103.405 184.675 ;
        RECT 103.925 184.385 104.205 184.845 ;
        RECT 104.395 184.385 104.795 185.185 ;
        RECT 104.965 185.915 105.920 186.135 ;
        RECT 106.780 186.135 107.065 186.595 ;
        RECT 107.235 186.305 107.505 186.765 ;
        RECT 106.780 185.915 107.735 186.135 ;
        RECT 104.965 185.015 105.175 185.915 ;
        RECT 105.345 185.185 106.035 185.745 ;
        RECT 106.665 185.185 107.355 185.745 ;
        RECT 107.525 185.015 107.735 185.915 ;
        RECT 104.965 184.845 105.920 185.015 ;
        RECT 105.195 184.215 105.465 184.675 ;
        RECT 105.635 184.385 105.920 184.845 ;
        RECT 106.780 184.845 107.735 185.015 ;
        RECT 107.905 185.745 108.305 186.595 ;
        RECT 108.495 186.135 108.775 186.595 ;
        RECT 109.295 186.305 109.620 186.765 ;
        RECT 108.495 185.915 109.620 186.135 ;
        RECT 107.905 185.185 109.000 185.745 ;
        RECT 109.170 185.455 109.620 185.915 ;
        RECT 109.790 185.625 110.175 186.595 ;
        RECT 110.460 186.135 110.745 186.595 ;
        RECT 110.915 186.305 111.185 186.765 ;
        RECT 110.460 185.915 111.415 186.135 ;
        RECT 106.780 184.385 107.065 184.845 ;
        RECT 107.235 184.215 107.505 184.675 ;
        RECT 107.905 184.385 108.305 185.185 ;
        RECT 109.170 185.125 109.725 185.455 ;
        RECT 109.170 185.015 109.620 185.125 ;
        RECT 108.495 184.845 109.620 185.015 ;
        RECT 109.895 184.955 110.175 185.625 ;
        RECT 110.345 185.185 111.035 185.745 ;
        RECT 111.205 185.015 111.415 185.915 ;
        RECT 108.495 184.385 108.775 184.845 ;
        RECT 109.295 184.215 109.620 184.675 ;
        RECT 109.790 184.385 110.175 184.955 ;
        RECT 110.460 184.845 111.415 185.015 ;
        RECT 111.585 185.745 111.985 186.595 ;
        RECT 112.175 186.135 112.455 186.595 ;
        RECT 112.975 186.305 113.300 186.765 ;
        RECT 112.175 185.915 113.300 186.135 ;
        RECT 111.585 185.185 112.680 185.745 ;
        RECT 112.850 185.455 113.300 185.915 ;
        RECT 113.470 185.625 113.855 186.595 ;
        RECT 110.460 184.385 110.745 184.845 ;
        RECT 110.915 184.215 111.185 184.675 ;
        RECT 111.585 184.385 111.985 185.185 ;
        RECT 112.850 185.125 113.405 185.455 ;
        RECT 112.850 185.015 113.300 185.125 ;
        RECT 112.175 184.845 113.300 185.015 ;
        RECT 113.575 184.955 113.855 185.625 ;
        RECT 114.025 185.675 115.235 186.765 ;
        RECT 115.410 186.330 120.755 186.765 ;
        RECT 120.930 186.330 126.275 186.765 ;
        RECT 114.025 185.135 114.545 185.675 ;
        RECT 114.715 184.965 115.235 185.505 ;
        RECT 117.000 185.080 117.350 186.330 ;
        RECT 112.175 184.385 112.455 184.845 ;
        RECT 112.975 184.215 113.300 184.675 ;
        RECT 113.470 184.385 113.855 184.955 ;
        RECT 114.025 184.215 115.235 184.965 ;
        RECT 118.830 184.760 119.170 185.590 ;
        RECT 122.520 185.080 122.870 186.330 ;
        RECT 126.445 185.675 127.655 186.765 ;
        RECT 124.350 184.760 124.690 185.590 ;
        RECT 126.445 185.135 126.965 185.675 ;
        RECT 127.135 184.965 127.655 185.505 ;
        RECT 115.410 184.215 120.755 184.760 ;
        RECT 120.930 184.215 126.275 184.760 ;
        RECT 126.445 184.215 127.655 184.965 ;
        RECT 14.580 184.045 127.740 184.215 ;
        RECT 14.665 183.295 15.875 184.045 ;
        RECT 16.510 183.500 21.855 184.045 ;
        RECT 14.665 182.755 15.185 183.295 ;
        RECT 15.355 182.585 15.875 183.125 ;
        RECT 14.665 181.495 15.875 182.585 ;
        RECT 18.100 181.930 18.450 183.180 ;
        RECT 19.930 182.670 20.270 183.500 ;
        RECT 22.115 183.495 22.285 183.875 ;
        RECT 22.465 183.665 22.795 184.045 ;
        RECT 22.115 183.325 22.780 183.495 ;
        RECT 22.975 183.370 23.235 183.875 ;
        RECT 22.045 182.775 22.375 183.145 ;
        RECT 22.610 183.070 22.780 183.325 ;
        RECT 22.610 182.740 22.895 183.070 ;
        RECT 22.610 182.595 22.780 182.740 ;
        RECT 22.115 182.425 22.780 182.595 ;
        RECT 23.065 182.570 23.235 183.370 ;
        RECT 16.510 181.495 21.855 181.930 ;
        RECT 22.115 181.665 22.285 182.425 ;
        RECT 22.465 181.495 22.795 182.255 ;
        RECT 22.965 181.665 23.235 182.570 ;
        RECT 23.405 183.305 23.790 183.875 ;
        RECT 23.960 183.585 24.285 184.045 ;
        RECT 24.805 183.415 25.085 183.875 ;
        RECT 23.405 182.635 23.685 183.305 ;
        RECT 23.960 183.245 25.085 183.415 ;
        RECT 23.960 183.135 24.410 183.245 ;
        RECT 23.855 182.805 24.410 183.135 ;
        RECT 25.275 183.075 25.675 183.875 ;
        RECT 26.075 183.585 26.345 184.045 ;
        RECT 26.515 183.415 26.800 183.875 ;
        RECT 23.405 181.665 23.790 182.635 ;
        RECT 23.960 182.345 24.410 182.805 ;
        RECT 24.580 182.515 25.675 183.075 ;
        RECT 23.960 182.125 25.085 182.345 ;
        RECT 23.960 181.495 24.285 181.955 ;
        RECT 24.805 181.665 25.085 182.125 ;
        RECT 25.275 181.665 25.675 182.515 ;
        RECT 25.845 183.245 26.800 183.415 ;
        RECT 27.200 183.415 27.485 183.875 ;
        RECT 27.655 183.585 27.925 184.045 ;
        RECT 27.200 183.245 28.155 183.415 ;
        RECT 25.845 182.345 26.055 183.245 ;
        RECT 26.225 182.515 26.915 183.075 ;
        RECT 27.085 182.515 27.775 183.075 ;
        RECT 27.945 182.345 28.155 183.245 ;
        RECT 25.845 182.125 26.800 182.345 ;
        RECT 26.075 181.495 26.345 181.955 ;
        RECT 26.515 181.665 26.800 182.125 ;
        RECT 27.200 182.125 28.155 182.345 ;
        RECT 28.325 183.075 28.725 183.875 ;
        RECT 28.915 183.415 29.195 183.875 ;
        RECT 29.715 183.585 30.040 184.045 ;
        RECT 28.915 183.245 30.040 183.415 ;
        RECT 30.210 183.305 30.595 183.875 ;
        RECT 29.590 183.135 30.040 183.245 ;
        RECT 28.325 182.515 29.420 183.075 ;
        RECT 29.590 182.805 30.145 183.135 ;
        RECT 27.200 181.665 27.485 182.125 ;
        RECT 27.655 181.495 27.925 181.955 ;
        RECT 28.325 181.665 28.725 182.515 ;
        RECT 29.590 182.345 30.040 182.805 ;
        RECT 30.315 182.635 30.595 183.305 ;
        RECT 28.915 182.125 30.040 182.345 ;
        RECT 28.915 181.665 29.195 182.125 ;
        RECT 29.715 181.495 30.040 181.955 ;
        RECT 30.210 181.665 30.595 182.635 ;
        RECT 30.770 183.305 31.025 183.875 ;
        RECT 31.195 183.645 31.525 184.045 ;
        RECT 31.950 183.510 32.480 183.875 ;
        RECT 31.950 183.475 32.125 183.510 ;
        RECT 31.195 183.305 32.125 183.475 ;
        RECT 32.670 183.365 32.945 183.875 ;
        RECT 30.770 182.635 30.940 183.305 ;
        RECT 31.195 183.135 31.365 183.305 ;
        RECT 31.110 182.805 31.365 183.135 ;
        RECT 31.590 182.805 31.785 183.135 ;
        RECT 30.770 181.665 31.105 182.635 ;
        RECT 31.275 181.495 31.445 182.635 ;
        RECT 31.615 181.835 31.785 182.805 ;
        RECT 31.955 182.175 32.125 183.305 ;
        RECT 32.295 182.515 32.465 183.315 ;
        RECT 32.665 183.195 32.945 183.365 ;
        RECT 32.670 182.715 32.945 183.195 ;
        RECT 33.115 182.515 33.305 183.875 ;
        RECT 33.485 183.510 33.995 184.045 ;
        RECT 34.215 183.235 34.460 183.840 ;
        RECT 35.365 183.275 37.035 184.045 ;
        RECT 37.205 183.320 37.495 184.045 ;
        RECT 37.780 183.415 38.065 183.875 ;
        RECT 38.235 183.585 38.505 184.045 ;
        RECT 33.505 183.065 34.735 183.235 ;
        RECT 32.295 182.345 33.305 182.515 ;
        RECT 33.475 182.500 34.225 182.690 ;
        RECT 31.955 182.005 33.080 182.175 ;
        RECT 33.475 181.835 33.645 182.500 ;
        RECT 34.395 182.255 34.735 183.065 ;
        RECT 31.615 181.665 33.645 181.835 ;
        RECT 33.815 181.495 33.985 182.255 ;
        RECT 34.220 181.845 34.735 182.255 ;
        RECT 35.365 182.585 36.115 183.105 ;
        RECT 36.285 182.755 37.035 183.275 ;
        RECT 37.780 183.245 38.735 183.415 ;
        RECT 35.365 181.495 37.035 182.585 ;
        RECT 37.205 181.495 37.495 182.660 ;
        RECT 37.665 182.515 38.355 183.075 ;
        RECT 38.525 182.345 38.735 183.245 ;
        RECT 37.780 182.125 38.735 182.345 ;
        RECT 38.905 183.075 39.305 183.875 ;
        RECT 39.495 183.415 39.775 183.875 ;
        RECT 40.295 183.585 40.620 184.045 ;
        RECT 39.495 183.245 40.620 183.415 ;
        RECT 40.790 183.305 41.175 183.875 ;
        RECT 40.170 183.135 40.620 183.245 ;
        RECT 38.905 182.515 40.000 183.075 ;
        RECT 40.170 182.805 40.725 183.135 ;
        RECT 37.780 181.665 38.065 182.125 ;
        RECT 38.235 181.495 38.505 181.955 ;
        RECT 38.905 181.665 39.305 182.515 ;
        RECT 40.170 182.345 40.620 182.805 ;
        RECT 40.895 182.635 41.175 183.305 ;
        RECT 41.460 183.415 41.745 183.875 ;
        RECT 41.915 183.585 42.185 184.045 ;
        RECT 41.460 183.245 42.415 183.415 ;
        RECT 39.495 182.125 40.620 182.345 ;
        RECT 39.495 181.665 39.775 182.125 ;
        RECT 40.295 181.495 40.620 181.955 ;
        RECT 40.790 181.665 41.175 182.635 ;
        RECT 41.345 182.515 42.035 183.075 ;
        RECT 42.205 182.345 42.415 183.245 ;
        RECT 41.460 182.125 42.415 182.345 ;
        RECT 42.585 183.075 42.985 183.875 ;
        RECT 43.175 183.415 43.455 183.875 ;
        RECT 43.975 183.585 44.300 184.045 ;
        RECT 43.175 183.245 44.300 183.415 ;
        RECT 44.470 183.305 44.855 183.875 ;
        RECT 43.850 183.135 44.300 183.245 ;
        RECT 42.585 182.515 43.680 183.075 ;
        RECT 43.850 182.805 44.405 183.135 ;
        RECT 41.460 181.665 41.745 182.125 ;
        RECT 41.915 181.495 42.185 181.955 ;
        RECT 42.585 181.665 42.985 182.515 ;
        RECT 43.850 182.345 44.300 182.805 ;
        RECT 44.575 182.635 44.855 183.305 ;
        RECT 45.140 183.415 45.425 183.875 ;
        RECT 45.595 183.585 45.865 184.045 ;
        RECT 45.140 183.245 46.095 183.415 ;
        RECT 43.175 182.125 44.300 182.345 ;
        RECT 43.175 181.665 43.455 182.125 ;
        RECT 43.975 181.495 44.300 181.955 ;
        RECT 44.470 181.665 44.855 182.635 ;
        RECT 45.025 182.515 45.715 183.075 ;
        RECT 45.885 182.345 46.095 183.245 ;
        RECT 45.140 182.125 46.095 182.345 ;
        RECT 46.265 183.075 46.665 183.875 ;
        RECT 46.855 183.415 47.135 183.875 ;
        RECT 47.655 183.585 47.980 184.045 ;
        RECT 46.855 183.245 47.980 183.415 ;
        RECT 48.150 183.305 48.535 183.875 ;
        RECT 47.530 183.135 47.980 183.245 ;
        RECT 46.265 182.515 47.360 183.075 ;
        RECT 47.530 182.805 48.085 183.135 ;
        RECT 45.140 181.665 45.425 182.125 ;
        RECT 45.595 181.495 45.865 181.955 ;
        RECT 46.265 181.665 46.665 182.515 ;
        RECT 47.530 182.345 47.980 182.805 ;
        RECT 48.255 182.635 48.535 183.305 ;
        RECT 46.855 182.125 47.980 182.345 ;
        RECT 46.855 181.665 47.135 182.125 ;
        RECT 47.655 181.495 47.980 181.955 ;
        RECT 48.150 181.665 48.535 182.635 ;
        RECT 48.705 183.370 48.965 183.875 ;
        RECT 49.145 183.665 49.475 184.045 ;
        RECT 49.655 183.495 49.825 183.875 ;
        RECT 48.705 182.570 48.875 183.370 ;
        RECT 49.160 183.325 49.825 183.495 ;
        RECT 50.085 183.370 50.345 183.875 ;
        RECT 50.525 183.665 50.855 184.045 ;
        RECT 51.035 183.495 51.205 183.875 ;
        RECT 49.160 183.070 49.330 183.325 ;
        RECT 49.045 182.740 49.330 183.070 ;
        RECT 49.565 182.775 49.895 183.145 ;
        RECT 49.160 182.595 49.330 182.740 ;
        RECT 48.705 181.665 48.975 182.570 ;
        RECT 49.160 182.425 49.825 182.595 ;
        RECT 49.145 181.495 49.475 182.255 ;
        RECT 49.655 181.665 49.825 182.425 ;
        RECT 50.085 182.570 50.255 183.370 ;
        RECT 50.540 183.325 51.205 183.495 ;
        RECT 51.555 183.495 51.725 183.875 ;
        RECT 51.905 183.665 52.235 184.045 ;
        RECT 51.555 183.325 52.220 183.495 ;
        RECT 52.415 183.370 52.675 183.875 ;
        RECT 52.945 183.580 53.195 184.045 ;
        RECT 53.365 183.405 53.535 183.875 ;
        RECT 53.785 183.585 53.955 184.045 ;
        RECT 54.205 183.405 54.375 183.875 ;
        RECT 54.625 183.585 54.795 184.045 ;
        RECT 55.045 183.405 55.215 183.875 ;
        RECT 55.585 183.585 55.850 184.045 ;
        RECT 50.540 183.070 50.710 183.325 ;
        RECT 50.425 182.740 50.710 183.070 ;
        RECT 50.945 182.775 51.275 183.145 ;
        RECT 51.485 182.775 51.815 183.145 ;
        RECT 52.050 183.070 52.220 183.325 ;
        RECT 50.540 182.595 50.710 182.740 ;
        RECT 52.050 182.740 52.335 183.070 ;
        RECT 52.050 182.595 52.220 182.740 ;
        RECT 50.085 181.665 50.355 182.570 ;
        RECT 50.540 182.425 51.205 182.595 ;
        RECT 50.525 181.495 50.855 182.255 ;
        RECT 51.035 181.665 51.205 182.425 ;
        RECT 51.555 182.425 52.220 182.595 ;
        RECT 52.505 182.570 52.675 183.370 ;
        RECT 51.555 181.665 51.725 182.425 ;
        RECT 51.905 181.495 52.235 182.255 ;
        RECT 52.405 181.665 52.675 182.570 ;
        RECT 52.845 183.225 55.215 183.405 ;
        RECT 56.525 183.275 59.115 184.045 ;
        RECT 52.845 182.635 53.195 183.225 ;
        RECT 53.365 182.805 55.875 183.055 ;
        RECT 52.845 182.465 55.295 182.635 ;
        RECT 52.845 182.445 53.615 182.465 ;
        RECT 52.945 181.495 53.115 181.955 ;
        RECT 53.285 181.665 53.615 182.445 ;
        RECT 53.785 181.495 53.955 182.295 ;
        RECT 54.125 181.665 54.455 182.465 ;
        RECT 54.625 181.495 54.795 182.295 ;
        RECT 54.965 181.665 55.295 182.465 ;
        RECT 55.555 181.495 55.850 182.635 ;
        RECT 56.525 182.585 57.735 183.105 ;
        RECT 57.905 182.755 59.115 183.275 ;
        RECT 59.345 183.225 59.555 184.045 ;
        RECT 59.725 183.245 60.055 183.875 ;
        RECT 59.725 182.645 59.975 183.245 ;
        RECT 60.225 183.225 60.455 184.045 ;
        RECT 61.125 183.275 62.795 184.045 ;
        RECT 62.965 183.320 63.255 184.045 ;
        RECT 63.885 183.275 66.475 184.045 ;
        RECT 66.915 183.650 67.245 184.045 ;
        RECT 67.415 183.475 67.615 183.830 ;
        RECT 67.785 183.645 68.115 184.045 ;
        RECT 68.285 183.475 68.485 183.820 ;
        RECT 60.145 182.805 60.475 183.055 ;
        RECT 56.525 181.495 59.115 182.585 ;
        RECT 59.345 181.495 59.555 182.635 ;
        RECT 59.725 181.665 60.055 182.645 ;
        RECT 60.225 181.495 60.455 182.635 ;
        RECT 61.125 182.585 61.875 183.105 ;
        RECT 62.045 182.755 62.795 183.275 ;
        RECT 61.125 181.495 62.795 182.585 ;
        RECT 62.965 181.495 63.255 182.660 ;
        RECT 63.885 182.585 65.095 183.105 ;
        RECT 65.265 182.755 66.475 183.275 ;
        RECT 66.645 183.305 68.485 183.475 ;
        RECT 68.655 183.305 68.985 184.045 ;
        RECT 69.220 183.475 69.390 183.725 ;
        RECT 69.220 183.305 69.695 183.475 ;
        RECT 63.885 181.495 66.475 182.585 ;
        RECT 66.645 181.680 66.905 183.305 ;
        RECT 67.085 182.335 67.305 183.135 ;
        RECT 67.545 182.515 67.845 183.135 ;
        RECT 68.015 182.515 68.345 183.135 ;
        RECT 68.515 182.515 68.835 183.135 ;
        RECT 69.005 182.515 69.355 183.135 ;
        RECT 69.525 182.335 69.695 183.305 ;
        RECT 69.865 183.225 70.125 184.045 ;
        RECT 70.295 183.405 70.625 183.875 ;
        RECT 70.795 183.575 70.965 184.045 ;
        RECT 71.135 183.405 71.465 183.875 ;
        RECT 71.635 183.575 72.360 184.045 ;
        RECT 72.530 183.405 72.860 183.875 ;
        RECT 73.030 183.575 73.200 184.045 ;
        RECT 73.370 183.405 73.700 183.875 ;
        RECT 70.295 183.225 73.700 183.405 ;
        RECT 73.870 183.235 74.075 184.045 ;
        RECT 73.495 183.055 73.700 183.225 ;
        RECT 74.245 183.225 74.600 183.750 ;
        RECT 74.770 183.305 75.020 184.045 ;
        RECT 75.690 183.475 75.860 183.725 ;
        RECT 75.385 183.305 75.860 183.475 ;
        RECT 76.095 183.305 76.425 184.045 ;
        RECT 76.595 183.475 76.795 183.820 ;
        RECT 76.965 183.645 77.295 184.045 ;
        RECT 77.465 183.475 77.665 183.830 ;
        RECT 77.835 183.650 78.165 184.045 ;
        RECT 76.595 183.305 78.435 183.475 ;
        RECT 74.245 183.055 74.415 183.225 ;
        RECT 69.880 182.845 71.020 183.055 ;
        RECT 71.200 182.845 72.415 183.055 ;
        RECT 72.595 182.845 73.315 183.055 ;
        RECT 73.495 182.675 73.815 183.055 ;
        RECT 74.100 182.885 74.415 183.055 ;
        RECT 67.085 182.125 69.695 182.335 ;
        RECT 69.865 182.505 71.885 182.675 ;
        RECT 68.655 181.495 68.985 181.945 ;
        RECT 69.865 181.665 70.205 182.505 ;
        RECT 70.375 181.495 70.585 182.335 ;
        RECT 70.755 181.665 71.005 182.505 ;
        RECT 71.175 181.835 71.385 182.335 ;
        RECT 71.555 182.005 71.885 182.505 ;
        RECT 72.055 182.505 73.240 182.675 ;
        RECT 72.055 182.005 72.440 182.505 ;
        RECT 72.610 181.835 72.820 182.335 ;
        RECT 71.175 181.665 72.820 181.835 ;
        RECT 72.990 181.835 73.240 182.505 ;
        RECT 73.410 182.505 73.815 182.675 ;
        RECT 73.410 182.005 73.660 182.505 ;
        RECT 73.830 181.835 74.075 182.335 ;
        RECT 72.990 181.665 74.075 181.835 ;
        RECT 74.245 182.095 74.415 182.885 ;
        RECT 74.585 182.845 75.215 183.055 ;
        RECT 74.965 182.175 75.215 182.845 ;
        RECT 75.385 182.335 75.555 183.305 ;
        RECT 75.725 182.515 76.075 183.135 ;
        RECT 76.245 182.515 76.565 183.135 ;
        RECT 76.735 182.515 77.065 183.135 ;
        RECT 77.235 182.515 77.535 183.135 ;
        RECT 77.775 182.335 77.995 183.135 ;
        RECT 75.385 182.125 77.995 182.335 ;
        RECT 74.245 181.680 74.600 182.095 ;
        RECT 74.770 181.495 75.020 181.995 ;
        RECT 76.095 181.495 76.425 181.945 ;
        RECT 78.175 181.680 78.435 183.305 ;
        RECT 79.530 183.335 79.785 183.865 ;
        RECT 79.955 183.585 80.260 184.045 ;
        RECT 80.505 183.665 81.575 183.835 ;
        RECT 79.530 182.685 79.740 183.335 ;
        RECT 80.505 183.310 80.825 183.665 ;
        RECT 80.500 183.135 80.825 183.310 ;
        RECT 79.910 182.835 80.825 183.135 ;
        RECT 80.995 183.095 81.235 183.495 ;
        RECT 81.405 183.435 81.575 183.665 ;
        RECT 81.745 183.605 81.935 184.045 ;
        RECT 82.105 183.595 83.055 183.875 ;
        RECT 83.275 183.685 83.625 183.855 ;
        RECT 81.405 183.265 81.935 183.435 ;
        RECT 79.910 182.805 80.650 182.835 ;
        RECT 79.530 181.805 79.785 182.685 ;
        RECT 79.955 181.495 80.260 182.635 ;
        RECT 80.480 182.215 80.650 182.805 ;
        RECT 80.995 182.725 81.535 183.095 ;
        RECT 81.715 182.985 81.935 183.265 ;
        RECT 82.105 182.815 82.275 183.595 ;
        RECT 81.870 182.645 82.275 182.815 ;
        RECT 82.445 182.805 82.795 183.425 ;
        RECT 81.870 182.555 82.040 182.645 ;
        RECT 82.965 182.635 83.175 183.425 ;
        RECT 80.820 182.385 82.040 182.555 ;
        RECT 82.500 182.475 83.175 182.635 ;
        RECT 80.480 182.045 81.280 182.215 ;
        RECT 80.600 181.495 80.930 181.875 ;
        RECT 81.110 181.755 81.280 182.045 ;
        RECT 81.870 182.005 82.040 182.385 ;
        RECT 82.210 182.465 83.175 182.475 ;
        RECT 83.365 183.295 83.625 183.685 ;
        RECT 83.835 183.585 84.165 184.045 ;
        RECT 85.040 183.655 85.895 183.825 ;
        RECT 86.100 183.655 86.595 183.825 ;
        RECT 86.765 183.685 87.095 184.045 ;
        RECT 83.365 182.605 83.535 183.295 ;
        RECT 83.705 182.945 83.875 183.125 ;
        RECT 84.045 183.115 84.835 183.365 ;
        RECT 85.040 182.945 85.210 183.655 ;
        RECT 85.380 183.145 85.735 183.365 ;
        RECT 83.705 182.775 85.395 182.945 ;
        RECT 82.210 182.175 82.670 182.465 ;
        RECT 83.365 182.435 84.865 182.605 ;
        RECT 83.365 182.295 83.535 182.435 ;
        RECT 82.975 182.125 83.535 182.295 ;
        RECT 81.450 181.495 81.700 181.955 ;
        RECT 81.870 181.665 82.740 182.005 ;
        RECT 82.975 181.665 83.145 182.125 ;
        RECT 83.980 182.095 85.055 182.265 ;
        RECT 83.315 181.495 83.685 181.955 ;
        RECT 83.980 181.755 84.150 182.095 ;
        RECT 84.320 181.495 84.650 181.925 ;
        RECT 84.885 181.755 85.055 182.095 ;
        RECT 85.225 181.995 85.395 182.775 ;
        RECT 85.565 182.555 85.735 183.145 ;
        RECT 85.905 182.745 86.255 183.365 ;
        RECT 85.565 182.165 86.030 182.555 ;
        RECT 86.425 182.295 86.595 183.655 ;
        RECT 86.765 182.465 87.225 183.515 ;
        RECT 86.200 182.125 86.595 182.295 ;
        RECT 86.200 181.995 86.370 182.125 ;
        RECT 85.225 181.665 85.905 181.995 ;
        RECT 86.120 181.665 86.370 181.995 ;
        RECT 86.540 181.495 86.790 181.955 ;
        RECT 86.960 181.680 87.285 182.465 ;
        RECT 87.455 181.665 87.625 183.785 ;
        RECT 87.795 183.665 88.125 184.045 ;
        RECT 88.295 183.495 88.550 183.785 ;
        RECT 87.800 183.325 88.550 183.495 ;
        RECT 87.800 182.335 88.030 183.325 ;
        RECT 88.725 183.320 89.015 184.045 ;
        RECT 89.245 183.225 89.455 184.045 ;
        RECT 89.625 183.245 89.955 183.875 ;
        RECT 88.200 182.505 88.550 183.155 ;
        RECT 87.800 182.165 88.550 182.335 ;
        RECT 87.795 181.495 88.125 181.995 ;
        RECT 88.295 181.665 88.550 182.165 ;
        RECT 88.725 181.495 89.015 182.660 ;
        RECT 89.625 182.645 89.875 183.245 ;
        RECT 90.125 183.225 90.355 184.045 ;
        RECT 90.565 183.295 91.775 184.045 ;
        RECT 90.045 182.805 90.375 183.055 ;
        RECT 89.245 181.495 89.455 182.635 ;
        RECT 89.625 181.665 89.955 182.645 ;
        RECT 90.125 181.495 90.355 182.635 ;
        RECT 90.565 182.585 91.085 183.125 ;
        RECT 91.255 182.755 91.775 183.295 ;
        RECT 91.945 183.275 95.455 184.045 ;
        RECT 91.945 182.585 93.635 183.105 ;
        RECT 93.805 182.755 95.455 183.275 ;
        RECT 95.900 183.235 96.145 183.840 ;
        RECT 96.365 183.510 96.875 184.045 ;
        RECT 95.625 183.065 96.855 183.235 ;
        RECT 90.565 181.495 91.775 182.585 ;
        RECT 91.945 181.495 95.455 182.585 ;
        RECT 95.625 182.255 95.965 183.065 ;
        RECT 96.135 182.500 96.885 182.690 ;
        RECT 95.625 181.845 96.140 182.255 ;
        RECT 96.375 181.495 96.545 182.255 ;
        RECT 96.715 181.835 96.885 182.500 ;
        RECT 97.055 182.515 97.245 183.875 ;
        RECT 97.415 183.705 97.690 183.875 ;
        RECT 97.415 183.535 97.695 183.705 ;
        RECT 97.415 182.715 97.690 183.535 ;
        RECT 97.880 183.510 98.410 183.875 ;
        RECT 98.835 183.645 99.165 184.045 ;
        RECT 98.235 183.475 98.410 183.510 ;
        RECT 97.895 182.515 98.065 183.315 ;
        RECT 97.055 182.345 98.065 182.515 ;
        RECT 98.235 183.305 99.165 183.475 ;
        RECT 99.335 183.305 99.590 183.875 ;
        RECT 98.235 182.175 98.405 183.305 ;
        RECT 98.995 183.135 99.165 183.305 ;
        RECT 97.280 182.005 98.405 182.175 ;
        RECT 98.575 182.805 98.770 183.135 ;
        RECT 98.995 182.805 99.250 183.135 ;
        RECT 98.575 181.835 98.745 182.805 ;
        RECT 99.420 182.635 99.590 183.305 ;
        RECT 99.765 183.275 102.355 184.045 ;
        RECT 96.715 181.665 98.745 181.835 ;
        RECT 98.915 181.495 99.085 182.635 ;
        RECT 99.255 181.665 99.590 182.635 ;
        RECT 99.765 182.585 100.975 183.105 ;
        RECT 101.145 182.755 102.355 183.275 ;
        RECT 102.800 183.235 103.045 183.840 ;
        RECT 103.265 183.510 103.775 184.045 ;
        RECT 102.525 183.065 103.755 183.235 ;
        RECT 99.765 181.495 102.355 182.585 ;
        RECT 102.525 182.255 102.865 183.065 ;
        RECT 103.035 182.500 103.785 182.690 ;
        RECT 102.525 181.845 103.040 182.255 ;
        RECT 103.275 181.495 103.445 182.255 ;
        RECT 103.615 181.835 103.785 182.500 ;
        RECT 103.955 182.515 104.145 183.875 ;
        RECT 104.315 183.365 104.590 183.875 ;
        RECT 104.780 183.510 105.310 183.875 ;
        RECT 105.735 183.645 106.065 184.045 ;
        RECT 105.135 183.475 105.310 183.510 ;
        RECT 104.315 183.195 104.595 183.365 ;
        RECT 104.315 182.715 104.590 183.195 ;
        RECT 104.795 182.515 104.965 183.315 ;
        RECT 103.955 182.345 104.965 182.515 ;
        RECT 105.135 183.305 106.065 183.475 ;
        RECT 106.235 183.305 106.490 183.875 ;
        RECT 105.135 182.175 105.305 183.305 ;
        RECT 105.895 183.135 106.065 183.305 ;
        RECT 104.180 182.005 105.305 182.175 ;
        RECT 105.475 182.805 105.670 183.135 ;
        RECT 105.895 182.805 106.150 183.135 ;
        RECT 105.475 181.835 105.645 182.805 ;
        RECT 106.320 182.635 106.490 183.305 ;
        RECT 103.615 181.665 105.645 181.835 ;
        RECT 105.815 181.495 105.985 182.635 ;
        RECT 106.155 181.665 106.490 182.635 ;
        RECT 106.665 183.245 107.005 183.875 ;
        RECT 107.175 183.245 107.425 184.045 ;
        RECT 107.615 183.395 107.945 183.875 ;
        RECT 108.115 183.585 108.340 184.045 ;
        RECT 108.510 183.395 108.840 183.875 ;
        RECT 106.665 182.685 106.840 183.245 ;
        RECT 107.615 183.225 108.840 183.395 ;
        RECT 109.470 183.265 109.970 183.875 ;
        RECT 107.010 182.885 107.705 183.055 ;
        RECT 106.665 182.635 106.895 182.685 ;
        RECT 107.535 182.635 107.705 182.885 ;
        RECT 107.880 182.855 108.300 183.055 ;
        RECT 108.470 182.855 108.800 183.055 ;
        RECT 108.970 182.855 109.300 183.055 ;
        RECT 109.470 182.635 109.640 183.265 ;
        RECT 110.620 183.235 110.865 183.840 ;
        RECT 111.085 183.510 111.595 184.045 ;
        RECT 110.345 183.065 111.575 183.235 ;
        RECT 109.825 182.805 110.175 183.055 ;
        RECT 106.665 181.665 107.005 182.635 ;
        RECT 107.175 181.495 107.345 182.635 ;
        RECT 107.535 182.465 109.970 182.635 ;
        RECT 107.615 181.495 107.865 182.295 ;
        RECT 108.510 181.665 108.840 182.465 ;
        RECT 109.140 181.495 109.470 182.295 ;
        RECT 109.640 181.665 109.970 182.465 ;
        RECT 110.345 182.255 110.685 183.065 ;
        RECT 110.855 182.500 111.605 182.690 ;
        RECT 110.345 181.845 110.860 182.255 ;
        RECT 111.095 181.495 111.265 182.255 ;
        RECT 111.435 181.835 111.605 182.500 ;
        RECT 111.775 182.515 111.965 183.875 ;
        RECT 112.135 183.025 112.410 183.875 ;
        RECT 112.600 183.510 113.130 183.875 ;
        RECT 113.555 183.645 113.885 184.045 ;
        RECT 112.955 183.475 113.130 183.510 ;
        RECT 112.135 182.855 112.415 183.025 ;
        RECT 112.135 182.715 112.410 182.855 ;
        RECT 112.615 182.515 112.785 183.315 ;
        RECT 111.775 182.345 112.785 182.515 ;
        RECT 112.955 183.305 113.885 183.475 ;
        RECT 114.055 183.305 114.310 183.875 ;
        RECT 114.485 183.320 114.775 184.045 ;
        RECT 115.870 183.335 116.125 183.865 ;
        RECT 116.295 183.585 116.600 184.045 ;
        RECT 116.845 183.665 117.915 183.835 ;
        RECT 112.955 182.175 113.125 183.305 ;
        RECT 113.715 183.135 113.885 183.305 ;
        RECT 112.000 182.005 113.125 182.175 ;
        RECT 113.295 182.805 113.490 183.135 ;
        RECT 113.715 182.805 113.970 183.135 ;
        RECT 113.295 181.835 113.465 182.805 ;
        RECT 114.140 182.635 114.310 183.305 ;
        RECT 115.870 182.685 116.080 183.335 ;
        RECT 116.845 183.310 117.165 183.665 ;
        RECT 116.840 183.135 117.165 183.310 ;
        RECT 116.250 182.835 117.165 183.135 ;
        RECT 117.335 183.095 117.575 183.495 ;
        RECT 117.745 183.435 117.915 183.665 ;
        RECT 118.085 183.605 118.275 184.045 ;
        RECT 118.445 183.595 119.395 183.875 ;
        RECT 119.615 183.685 119.965 183.855 ;
        RECT 117.745 183.265 118.275 183.435 ;
        RECT 116.250 182.805 116.990 182.835 ;
        RECT 111.435 181.665 113.465 181.835 ;
        RECT 113.635 181.495 113.805 182.635 ;
        RECT 113.975 181.665 114.310 182.635 ;
        RECT 114.485 181.495 114.775 182.660 ;
        RECT 115.870 181.805 116.125 182.685 ;
        RECT 116.295 181.495 116.600 182.635 ;
        RECT 116.820 182.215 116.990 182.805 ;
        RECT 117.335 182.725 117.875 183.095 ;
        RECT 118.055 182.985 118.275 183.265 ;
        RECT 118.445 182.815 118.615 183.595 ;
        RECT 118.210 182.645 118.615 182.815 ;
        RECT 118.785 182.805 119.135 183.425 ;
        RECT 118.210 182.555 118.380 182.645 ;
        RECT 119.305 182.635 119.515 183.425 ;
        RECT 117.160 182.385 118.380 182.555 ;
        RECT 118.840 182.475 119.515 182.635 ;
        RECT 116.820 182.045 117.620 182.215 ;
        RECT 116.940 181.495 117.270 181.875 ;
        RECT 117.450 181.755 117.620 182.045 ;
        RECT 118.210 182.005 118.380 182.385 ;
        RECT 118.550 182.465 119.515 182.475 ;
        RECT 119.705 183.295 119.965 183.685 ;
        RECT 120.175 183.585 120.505 184.045 ;
        RECT 121.380 183.655 122.235 183.825 ;
        RECT 122.440 183.655 122.935 183.825 ;
        RECT 123.105 183.685 123.435 184.045 ;
        RECT 119.705 182.605 119.875 183.295 ;
        RECT 120.045 182.945 120.215 183.125 ;
        RECT 120.385 183.115 121.175 183.365 ;
        RECT 121.380 182.945 121.550 183.655 ;
        RECT 121.720 183.145 122.075 183.365 ;
        RECT 120.045 182.775 121.735 182.945 ;
        RECT 118.550 182.175 119.010 182.465 ;
        RECT 119.705 182.435 121.205 182.605 ;
        RECT 119.705 182.295 119.875 182.435 ;
        RECT 119.315 182.125 119.875 182.295 ;
        RECT 117.790 181.495 118.040 181.955 ;
        RECT 118.210 181.665 119.080 182.005 ;
        RECT 119.315 181.665 119.485 182.125 ;
        RECT 120.320 182.095 121.395 182.265 ;
        RECT 119.655 181.495 120.025 181.955 ;
        RECT 120.320 181.755 120.490 182.095 ;
        RECT 120.660 181.495 120.990 181.925 ;
        RECT 121.225 181.755 121.395 182.095 ;
        RECT 121.565 181.995 121.735 182.775 ;
        RECT 121.905 182.555 122.075 183.145 ;
        RECT 122.245 182.745 122.595 183.365 ;
        RECT 121.905 182.165 122.370 182.555 ;
        RECT 122.765 182.295 122.935 183.655 ;
        RECT 123.105 182.465 123.565 183.515 ;
        RECT 122.540 182.125 122.935 182.295 ;
        RECT 122.540 181.995 122.710 182.125 ;
        RECT 121.565 181.665 122.245 181.995 ;
        RECT 122.460 181.665 122.710 181.995 ;
        RECT 122.880 181.495 123.130 181.955 ;
        RECT 123.300 181.680 123.625 182.465 ;
        RECT 123.795 181.665 123.965 183.785 ;
        RECT 124.135 183.665 124.465 184.045 ;
        RECT 124.635 183.495 124.890 183.785 ;
        RECT 124.140 183.325 124.890 183.495 ;
        RECT 124.140 182.335 124.370 183.325 ;
        RECT 125.065 183.295 126.275 184.045 ;
        RECT 126.445 183.295 127.655 184.045 ;
        RECT 124.540 182.505 124.890 183.155 ;
        RECT 125.065 182.585 125.585 183.125 ;
        RECT 125.755 182.755 126.275 183.295 ;
        RECT 126.445 182.585 126.965 183.125 ;
        RECT 127.135 182.755 127.655 183.295 ;
        RECT 124.140 182.165 124.890 182.335 ;
        RECT 124.135 181.495 124.465 181.995 ;
        RECT 124.635 181.665 124.890 182.165 ;
        RECT 125.065 181.495 126.275 182.585 ;
        RECT 126.445 181.495 127.655 182.585 ;
        RECT 14.580 181.325 127.740 181.495 ;
        RECT 14.665 180.235 15.875 181.325 ;
        RECT 14.665 179.525 15.185 180.065 ;
        RECT 15.355 179.695 15.875 180.235 ;
        RECT 16.045 180.235 18.635 181.325 ;
        RECT 18.810 180.890 24.155 181.325 ;
        RECT 16.045 179.715 17.255 180.235 ;
        RECT 17.425 179.545 18.635 180.065 ;
        RECT 20.400 179.640 20.750 180.890 ;
        RECT 24.325 180.160 24.615 181.325 ;
        RECT 24.790 180.655 25.045 181.155 ;
        RECT 25.215 180.825 25.545 181.325 ;
        RECT 24.790 180.485 25.540 180.655 ;
        RECT 14.665 178.775 15.875 179.525 ;
        RECT 16.045 178.775 18.635 179.545 ;
        RECT 22.230 179.320 22.570 180.150 ;
        RECT 24.790 179.665 25.140 180.315 ;
        RECT 18.810 178.775 24.155 179.320 ;
        RECT 24.325 178.775 24.615 179.500 ;
        RECT 25.310 179.495 25.540 180.485 ;
        RECT 24.790 179.325 25.540 179.495 ;
        RECT 24.790 179.035 25.045 179.325 ;
        RECT 25.215 178.775 25.545 179.155 ;
        RECT 25.715 179.035 25.885 181.155 ;
        RECT 26.055 180.355 26.380 181.140 ;
        RECT 26.550 180.865 26.800 181.325 ;
        RECT 26.970 180.825 27.220 181.155 ;
        RECT 27.435 180.825 28.115 181.155 ;
        RECT 26.970 180.695 27.140 180.825 ;
        RECT 26.745 180.525 27.140 180.695 ;
        RECT 26.115 179.305 26.575 180.355 ;
        RECT 26.745 179.165 26.915 180.525 ;
        RECT 27.310 180.265 27.775 180.655 ;
        RECT 27.085 179.455 27.435 180.075 ;
        RECT 27.605 179.675 27.775 180.265 ;
        RECT 27.945 180.045 28.115 180.825 ;
        RECT 28.285 180.725 28.455 181.065 ;
        RECT 28.690 180.895 29.020 181.325 ;
        RECT 29.190 180.725 29.360 181.065 ;
        RECT 29.655 180.865 30.025 181.325 ;
        RECT 28.285 180.555 29.360 180.725 ;
        RECT 30.195 180.695 30.365 181.155 ;
        RECT 30.600 180.815 31.470 181.155 ;
        RECT 31.640 180.865 31.890 181.325 ;
        RECT 29.805 180.525 30.365 180.695 ;
        RECT 29.805 180.385 29.975 180.525 ;
        RECT 28.475 180.215 29.975 180.385 ;
        RECT 30.670 180.355 31.130 180.645 ;
        RECT 27.945 179.875 29.635 180.045 ;
        RECT 27.605 179.455 27.960 179.675 ;
        RECT 28.130 179.165 28.300 179.875 ;
        RECT 28.505 179.455 29.295 179.705 ;
        RECT 29.465 179.695 29.635 179.875 ;
        RECT 29.805 179.525 29.975 180.215 ;
        RECT 26.245 178.775 26.575 179.135 ;
        RECT 26.745 178.995 27.240 179.165 ;
        RECT 27.445 178.995 28.300 179.165 ;
        RECT 29.175 178.775 29.505 179.235 ;
        RECT 29.715 179.135 29.975 179.525 ;
        RECT 30.165 180.345 31.130 180.355 ;
        RECT 31.300 180.435 31.470 180.815 ;
        RECT 32.060 180.775 32.230 181.065 ;
        RECT 32.410 180.945 32.740 181.325 ;
        RECT 32.060 180.605 32.860 180.775 ;
        RECT 30.165 180.185 30.840 180.345 ;
        RECT 31.300 180.265 32.520 180.435 ;
        RECT 30.165 179.395 30.375 180.185 ;
        RECT 31.300 180.175 31.470 180.265 ;
        RECT 30.545 179.395 30.895 180.015 ;
        RECT 31.065 180.005 31.470 180.175 ;
        RECT 31.065 179.225 31.235 180.005 ;
        RECT 31.405 179.555 31.625 179.835 ;
        RECT 31.805 179.725 32.345 180.095 ;
        RECT 32.690 180.015 32.860 180.605 ;
        RECT 33.080 180.185 33.385 181.325 ;
        RECT 33.555 180.135 33.810 181.015 ;
        RECT 32.690 179.985 33.430 180.015 ;
        RECT 31.405 179.385 31.935 179.555 ;
        RECT 29.715 178.965 30.065 179.135 ;
        RECT 30.285 178.945 31.235 179.225 ;
        RECT 31.405 178.775 31.595 179.215 ;
        RECT 31.765 179.155 31.935 179.385 ;
        RECT 32.105 179.325 32.345 179.725 ;
        RECT 32.515 179.685 33.430 179.985 ;
        RECT 32.515 179.510 32.840 179.685 ;
        RECT 32.515 179.155 32.835 179.510 ;
        RECT 33.600 179.485 33.810 180.135 ;
        RECT 31.765 178.985 32.835 179.155 ;
        RECT 33.080 178.775 33.385 179.235 ;
        RECT 33.555 178.955 33.810 179.485 ;
        RECT 33.985 180.185 34.370 181.155 ;
        RECT 34.540 180.865 34.865 181.325 ;
        RECT 35.385 180.695 35.665 181.155 ;
        RECT 34.540 180.475 35.665 180.695 ;
        RECT 33.985 179.515 34.265 180.185 ;
        RECT 34.540 180.015 34.990 180.475 ;
        RECT 35.855 180.305 36.255 181.155 ;
        RECT 36.655 180.865 36.925 181.325 ;
        RECT 37.095 180.695 37.380 181.155 ;
        RECT 34.435 179.685 34.990 180.015 ;
        RECT 35.160 179.745 36.255 180.305 ;
        RECT 34.540 179.575 34.990 179.685 ;
        RECT 33.985 178.945 34.370 179.515 ;
        RECT 34.540 179.405 35.665 179.575 ;
        RECT 34.540 178.775 34.865 179.235 ;
        RECT 35.385 178.945 35.665 179.405 ;
        RECT 35.855 178.945 36.255 179.745 ;
        RECT 36.425 180.475 37.380 180.695 ;
        RECT 36.425 179.575 36.635 180.475 ;
        RECT 36.805 179.745 37.495 180.305 ;
        RECT 38.125 180.185 38.465 181.155 ;
        RECT 38.635 180.185 38.805 181.325 ;
        RECT 39.075 180.525 39.325 181.325 ;
        RECT 39.970 180.355 40.300 181.155 ;
        RECT 40.600 180.525 40.930 181.325 ;
        RECT 41.100 180.355 41.430 181.155 ;
        RECT 38.995 180.185 41.430 180.355 ;
        RECT 42.265 180.185 42.605 181.155 ;
        RECT 42.775 180.185 42.945 181.325 ;
        RECT 43.215 180.525 43.465 181.325 ;
        RECT 44.110 180.355 44.440 181.155 ;
        RECT 44.740 180.525 45.070 181.325 ;
        RECT 45.240 180.355 45.570 181.155 ;
        RECT 43.135 180.185 45.570 180.355 ;
        RECT 45.945 180.565 46.460 180.975 ;
        RECT 46.695 180.565 46.865 181.325 ;
        RECT 47.035 180.985 49.065 181.155 ;
        RECT 38.125 179.625 38.300 180.185 ;
        RECT 38.995 179.935 39.165 180.185 ;
        RECT 38.470 179.765 39.165 179.935 ;
        RECT 39.340 179.765 39.760 179.965 ;
        RECT 39.930 179.765 40.260 179.965 ;
        RECT 40.430 179.765 40.760 179.965 ;
        RECT 38.125 179.575 38.355 179.625 ;
        RECT 36.425 179.405 37.380 179.575 ;
        RECT 36.655 178.775 36.925 179.235 ;
        RECT 37.095 178.945 37.380 179.405 ;
        RECT 38.125 178.945 38.465 179.575 ;
        RECT 38.635 178.775 38.885 179.575 ;
        RECT 39.075 179.425 40.300 179.595 ;
        RECT 39.075 178.945 39.405 179.425 ;
        RECT 39.575 178.775 39.800 179.235 ;
        RECT 39.970 178.945 40.300 179.425 ;
        RECT 40.930 179.555 41.100 180.185 ;
        RECT 41.285 179.765 41.635 180.015 ;
        RECT 42.265 179.575 42.440 180.185 ;
        RECT 43.135 179.935 43.305 180.185 ;
        RECT 42.610 179.765 43.305 179.935 ;
        RECT 43.480 179.765 43.900 179.965 ;
        RECT 44.070 179.765 44.400 179.965 ;
        RECT 44.570 179.765 44.900 179.965 ;
        RECT 40.930 178.945 41.430 179.555 ;
        RECT 42.265 178.945 42.605 179.575 ;
        RECT 42.775 178.775 43.025 179.575 ;
        RECT 43.215 179.425 44.440 179.595 ;
        RECT 43.215 178.945 43.545 179.425 ;
        RECT 43.715 178.775 43.940 179.235 ;
        RECT 44.110 178.945 44.440 179.425 ;
        RECT 45.070 179.555 45.240 180.185 ;
        RECT 45.425 179.765 45.775 180.015 ;
        RECT 45.945 179.755 46.285 180.565 ;
        RECT 47.035 180.320 47.205 180.985 ;
        RECT 47.600 180.645 48.725 180.815 ;
        RECT 46.455 180.130 47.205 180.320 ;
        RECT 47.375 180.305 48.385 180.475 ;
        RECT 45.945 179.585 47.175 179.755 ;
        RECT 45.070 178.945 45.570 179.555 ;
        RECT 46.220 178.980 46.465 179.585 ;
        RECT 46.685 178.775 47.195 179.310 ;
        RECT 47.375 178.945 47.565 180.305 ;
        RECT 47.735 179.285 48.010 180.105 ;
        RECT 48.215 179.505 48.385 180.305 ;
        RECT 48.555 179.515 48.725 180.645 ;
        RECT 48.895 180.015 49.065 180.985 ;
        RECT 49.235 180.185 49.405 181.325 ;
        RECT 49.575 180.185 49.910 181.155 ;
        RECT 48.895 179.685 49.090 180.015 ;
        RECT 49.315 179.685 49.570 180.015 ;
        RECT 49.315 179.515 49.485 179.685 ;
        RECT 49.740 179.515 49.910 180.185 ;
        RECT 50.085 180.160 50.375 181.325 ;
        RECT 50.660 180.695 50.945 181.155 ;
        RECT 51.115 180.865 51.385 181.325 ;
        RECT 50.660 180.475 51.615 180.695 ;
        RECT 50.545 179.745 51.235 180.305 ;
        RECT 51.405 179.575 51.615 180.475 ;
        RECT 48.555 179.345 49.485 179.515 ;
        RECT 48.555 179.310 48.730 179.345 ;
        RECT 47.735 179.115 48.015 179.285 ;
        RECT 47.735 178.945 48.010 179.115 ;
        RECT 48.200 178.945 48.730 179.310 ;
        RECT 49.155 178.775 49.485 179.175 ;
        RECT 49.655 178.945 49.910 179.515 ;
        RECT 50.085 178.775 50.375 179.500 ;
        RECT 50.660 179.405 51.615 179.575 ;
        RECT 51.785 180.305 52.185 181.155 ;
        RECT 52.375 180.695 52.655 181.155 ;
        RECT 53.175 180.865 53.500 181.325 ;
        RECT 52.375 180.475 53.500 180.695 ;
        RECT 51.785 179.745 52.880 180.305 ;
        RECT 53.050 180.015 53.500 180.475 ;
        RECT 53.670 180.185 54.055 181.155 ;
        RECT 50.660 178.945 50.945 179.405 ;
        RECT 51.115 178.775 51.385 179.235 ;
        RECT 51.785 178.945 52.185 179.745 ;
        RECT 53.050 179.685 53.605 180.015 ;
        RECT 53.050 179.575 53.500 179.685 ;
        RECT 52.375 179.405 53.500 179.575 ;
        RECT 53.775 179.515 54.055 180.185 ;
        RECT 54.225 180.235 55.895 181.325 ;
        RECT 54.225 179.715 54.975 180.235 ;
        RECT 56.070 180.185 56.405 181.155 ;
        RECT 56.575 180.185 56.745 181.325 ;
        RECT 56.915 180.985 58.945 181.155 ;
        RECT 55.145 179.545 55.895 180.065 ;
        RECT 52.375 178.945 52.655 179.405 ;
        RECT 53.175 178.775 53.500 179.235 ;
        RECT 53.670 178.945 54.055 179.515 ;
        RECT 54.225 178.775 55.895 179.545 ;
        RECT 56.070 179.515 56.240 180.185 ;
        RECT 56.915 180.015 57.085 180.985 ;
        RECT 56.410 179.685 56.665 180.015 ;
        RECT 56.890 179.685 57.085 180.015 ;
        RECT 57.255 180.645 58.380 180.815 ;
        RECT 56.495 179.515 56.665 179.685 ;
        RECT 57.255 179.515 57.425 180.645 ;
        RECT 56.070 178.945 56.325 179.515 ;
        RECT 56.495 179.345 57.425 179.515 ;
        RECT 57.595 180.305 58.605 180.475 ;
        RECT 57.595 179.505 57.765 180.305 ;
        RECT 57.250 179.310 57.425 179.345 ;
        RECT 56.495 178.775 56.825 179.175 ;
        RECT 57.250 178.945 57.780 179.310 ;
        RECT 57.970 179.285 58.245 180.105 ;
        RECT 57.965 179.115 58.245 179.285 ;
        RECT 57.970 178.945 58.245 179.115 ;
        RECT 58.415 178.945 58.605 180.305 ;
        RECT 58.775 180.320 58.945 180.985 ;
        RECT 59.115 180.565 59.285 181.325 ;
        RECT 59.520 180.565 60.035 180.975 ;
        RECT 58.775 180.130 59.525 180.320 ;
        RECT 59.695 179.755 60.035 180.565 ;
        RECT 60.260 180.455 60.545 181.325 ;
        RECT 60.715 180.695 60.975 181.155 ;
        RECT 61.150 180.865 61.405 181.325 ;
        RECT 61.575 180.695 61.835 181.155 ;
        RECT 60.715 180.525 61.835 180.695 ;
        RECT 62.005 180.525 62.315 181.325 ;
        RECT 60.715 180.275 60.975 180.525 ;
        RECT 62.485 180.355 62.795 181.155 ;
        RECT 58.805 179.585 60.035 179.755 ;
        RECT 60.220 180.105 60.975 180.275 ;
        RECT 61.765 180.185 62.795 180.355 ;
        RECT 60.220 179.595 60.625 180.105 ;
        RECT 61.765 179.935 61.935 180.185 ;
        RECT 60.795 179.765 61.935 179.935 ;
        RECT 58.785 178.775 59.295 179.310 ;
        RECT 59.515 178.980 59.760 179.585 ;
        RECT 60.220 179.425 61.870 179.595 ;
        RECT 62.105 179.445 62.455 180.015 ;
        RECT 60.265 178.775 60.545 179.255 ;
        RECT 60.715 179.035 60.975 179.425 ;
        RECT 61.150 178.775 61.405 179.255 ;
        RECT 61.575 179.035 61.870 179.425 ;
        RECT 62.625 179.275 62.795 180.185 ;
        RECT 62.965 180.235 65.555 181.325 ;
        RECT 62.965 179.715 64.175 180.235 ;
        RECT 65.765 180.185 65.995 181.325 ;
        RECT 66.165 180.175 66.495 181.155 ;
        RECT 66.665 180.185 66.875 181.325 ;
        RECT 67.110 180.175 67.370 181.325 ;
        RECT 67.545 180.250 67.800 181.155 ;
        RECT 67.970 180.565 68.300 181.325 ;
        RECT 68.515 180.395 68.685 181.155 ;
        RECT 64.345 179.545 65.555 180.065 ;
        RECT 65.745 179.765 66.075 180.015 ;
        RECT 62.050 178.775 62.325 179.255 ;
        RECT 62.495 178.945 62.795 179.275 ;
        RECT 62.965 178.775 65.555 179.545 ;
        RECT 65.765 178.775 65.995 179.595 ;
        RECT 66.245 179.575 66.495 180.175 ;
        RECT 66.165 178.945 66.495 179.575 ;
        RECT 66.665 178.775 66.875 179.595 ;
        RECT 67.110 178.775 67.370 179.615 ;
        RECT 67.545 179.520 67.715 180.250 ;
        RECT 67.970 180.225 68.685 180.395 ;
        RECT 68.945 180.355 69.255 181.155 ;
        RECT 69.425 180.525 69.735 181.325 ;
        RECT 69.905 180.695 70.165 181.155 ;
        RECT 70.335 180.865 70.590 181.325 ;
        RECT 70.765 180.695 71.025 181.155 ;
        RECT 69.905 180.525 71.025 180.695 ;
        RECT 67.970 180.015 68.140 180.225 ;
        RECT 68.945 180.185 69.975 180.355 ;
        RECT 67.885 179.685 68.140 180.015 ;
        RECT 67.545 178.945 67.800 179.520 ;
        RECT 67.970 179.495 68.140 179.685 ;
        RECT 68.420 179.675 68.775 180.045 ;
        RECT 67.970 179.325 68.685 179.495 ;
        RECT 67.970 178.775 68.300 179.155 ;
        RECT 68.515 178.945 68.685 179.325 ;
        RECT 68.945 179.275 69.115 180.185 ;
        RECT 69.285 179.445 69.635 180.015 ;
        RECT 69.805 179.935 69.975 180.185 ;
        RECT 70.765 180.275 71.025 180.525 ;
        RECT 71.195 180.455 71.480 181.325 ;
        RECT 70.765 180.105 71.520 180.275 ;
        RECT 69.805 179.765 70.945 179.935 ;
        RECT 71.115 179.595 71.520 180.105 ;
        RECT 69.870 179.425 71.520 179.595 ;
        RECT 71.705 179.515 71.965 181.140 ;
        RECT 73.715 180.875 74.045 181.325 ;
        RECT 72.145 180.485 74.755 180.695 ;
        RECT 72.145 179.685 72.365 180.485 ;
        RECT 72.605 179.685 72.905 180.305 ;
        RECT 73.075 179.685 73.405 180.305 ;
        RECT 73.575 179.685 73.895 180.305 ;
        RECT 74.065 179.685 74.415 180.305 ;
        RECT 74.585 179.515 74.755 180.485 ;
        RECT 75.845 180.160 76.135 181.325 ;
        RECT 76.420 180.695 76.705 181.155 ;
        RECT 76.875 180.865 77.145 181.325 ;
        RECT 76.420 180.475 77.375 180.695 ;
        RECT 76.305 179.745 76.995 180.305 ;
        RECT 77.165 179.575 77.375 180.475 ;
        RECT 68.945 178.945 69.245 179.275 ;
        RECT 69.415 178.775 69.690 179.255 ;
        RECT 69.870 179.035 70.165 179.425 ;
        RECT 70.335 178.775 70.590 179.255 ;
        RECT 70.765 179.035 71.025 179.425 ;
        RECT 71.705 179.345 73.545 179.515 ;
        RECT 71.195 178.775 71.475 179.255 ;
        RECT 71.975 178.775 72.305 179.170 ;
        RECT 72.475 178.990 72.675 179.345 ;
        RECT 72.845 178.775 73.175 179.175 ;
        RECT 73.345 179.000 73.545 179.345 ;
        RECT 73.715 178.775 74.045 179.515 ;
        RECT 74.280 179.345 74.755 179.515 ;
        RECT 74.280 179.095 74.450 179.345 ;
        RECT 75.845 178.775 76.135 179.500 ;
        RECT 76.420 179.405 77.375 179.575 ;
        RECT 77.545 180.305 77.945 181.155 ;
        RECT 78.135 180.695 78.415 181.155 ;
        RECT 78.935 180.865 79.260 181.325 ;
        RECT 78.135 180.475 79.260 180.695 ;
        RECT 77.545 179.745 78.640 180.305 ;
        RECT 78.810 180.015 79.260 180.475 ;
        RECT 79.430 180.185 79.815 181.155 ;
        RECT 80.190 180.355 80.520 181.155 ;
        RECT 80.690 180.525 81.020 181.325 ;
        RECT 81.320 180.355 81.650 181.155 ;
        RECT 82.295 180.525 82.545 181.325 ;
        RECT 80.190 180.185 82.625 180.355 ;
        RECT 82.815 180.185 82.985 181.325 ;
        RECT 83.155 180.185 83.495 181.155 ;
        RECT 76.420 178.945 76.705 179.405 ;
        RECT 76.875 178.775 77.145 179.235 ;
        RECT 77.545 178.945 77.945 179.745 ;
        RECT 78.810 179.685 79.365 180.015 ;
        RECT 78.810 179.575 79.260 179.685 ;
        RECT 78.135 179.405 79.260 179.575 ;
        RECT 79.535 179.515 79.815 180.185 ;
        RECT 79.985 179.765 80.335 180.015 ;
        RECT 80.520 179.555 80.690 180.185 ;
        RECT 80.860 179.765 81.190 179.965 ;
        RECT 81.360 179.765 81.690 179.965 ;
        RECT 81.860 179.765 82.280 179.965 ;
        RECT 82.455 179.935 82.625 180.185 ;
        RECT 82.455 179.765 83.150 179.935 ;
        RECT 78.135 178.945 78.415 179.405 ;
        RECT 78.935 178.775 79.260 179.235 ;
        RECT 79.430 178.945 79.815 179.515 ;
        RECT 80.190 178.945 80.690 179.555 ;
        RECT 81.320 179.425 82.545 179.595 ;
        RECT 83.320 179.575 83.495 180.185 ;
        RECT 83.665 180.235 85.335 181.325 ;
        RECT 85.505 180.565 86.020 180.975 ;
        RECT 86.255 180.565 86.425 181.325 ;
        RECT 86.595 180.985 88.625 181.155 ;
        RECT 83.665 179.715 84.415 180.235 ;
        RECT 81.320 178.945 81.650 179.425 ;
        RECT 81.820 178.775 82.045 179.235 ;
        RECT 82.215 178.945 82.545 179.425 ;
        RECT 82.735 178.775 82.985 179.575 ;
        RECT 83.155 178.945 83.495 179.575 ;
        RECT 84.585 179.545 85.335 180.065 ;
        RECT 85.505 179.755 85.845 180.565 ;
        RECT 86.595 180.320 86.765 180.985 ;
        RECT 87.160 180.645 88.285 180.815 ;
        RECT 86.015 180.130 86.765 180.320 ;
        RECT 86.935 180.305 87.945 180.475 ;
        RECT 85.505 179.585 86.735 179.755 ;
        RECT 83.665 178.775 85.335 179.545 ;
        RECT 85.780 178.980 86.025 179.585 ;
        RECT 86.245 178.775 86.755 179.310 ;
        RECT 86.935 178.945 87.125 180.305 ;
        RECT 87.295 179.285 87.570 180.105 ;
        RECT 87.775 179.505 87.945 180.305 ;
        RECT 88.115 179.515 88.285 180.645 ;
        RECT 88.455 180.015 88.625 180.985 ;
        RECT 88.795 180.185 88.965 181.325 ;
        RECT 89.135 180.185 89.470 181.155 ;
        RECT 88.455 179.685 88.650 180.015 ;
        RECT 88.875 179.685 89.130 180.015 ;
        RECT 88.875 179.515 89.045 179.685 ;
        RECT 89.300 179.515 89.470 180.185 ;
        RECT 88.115 179.345 89.045 179.515 ;
        RECT 88.115 179.310 88.290 179.345 ;
        RECT 87.295 179.115 87.575 179.285 ;
        RECT 87.295 178.945 87.570 179.115 ;
        RECT 87.760 178.945 88.290 179.310 ;
        RECT 88.715 178.775 89.045 179.175 ;
        RECT 89.215 178.945 89.470 179.515 ;
        RECT 89.645 180.250 89.915 181.155 ;
        RECT 90.085 180.565 90.415 181.325 ;
        RECT 90.595 180.395 90.765 181.155 ;
        RECT 89.645 179.450 89.815 180.250 ;
        RECT 90.100 180.225 90.765 180.395 ;
        RECT 90.100 180.080 90.270 180.225 ;
        RECT 91.065 180.185 91.295 181.325 ;
        RECT 91.465 180.175 91.795 181.155 ;
        RECT 91.965 180.185 92.175 181.325 ;
        RECT 89.985 179.750 90.270 180.080 ;
        RECT 90.100 179.495 90.270 179.750 ;
        RECT 90.505 179.675 90.835 180.045 ;
        RECT 91.045 179.765 91.375 180.015 ;
        RECT 89.645 178.945 89.905 179.450 ;
        RECT 90.100 179.325 90.765 179.495 ;
        RECT 90.085 178.775 90.415 179.155 ;
        RECT 90.595 178.945 90.765 179.325 ;
        RECT 91.065 178.775 91.295 179.595 ;
        RECT 91.545 179.575 91.795 180.175 ;
        RECT 92.410 180.135 92.665 181.015 ;
        RECT 92.835 180.185 93.140 181.325 ;
        RECT 93.480 180.945 93.810 181.325 ;
        RECT 93.990 180.775 94.160 181.065 ;
        RECT 94.330 180.865 94.580 181.325 ;
        RECT 93.360 180.605 94.160 180.775 ;
        RECT 94.750 180.815 95.620 181.155 ;
        RECT 91.465 178.945 91.795 179.575 ;
        RECT 91.965 178.775 92.175 179.595 ;
        RECT 92.410 179.485 92.620 180.135 ;
        RECT 93.360 180.015 93.530 180.605 ;
        RECT 94.750 180.435 94.920 180.815 ;
        RECT 95.855 180.695 96.025 181.155 ;
        RECT 96.195 180.865 96.565 181.325 ;
        RECT 96.860 180.725 97.030 181.065 ;
        RECT 97.200 180.895 97.530 181.325 ;
        RECT 97.765 180.725 97.935 181.065 ;
        RECT 93.700 180.265 94.920 180.435 ;
        RECT 95.090 180.355 95.550 180.645 ;
        RECT 95.855 180.525 96.415 180.695 ;
        RECT 96.860 180.555 97.935 180.725 ;
        RECT 98.105 180.825 98.785 181.155 ;
        RECT 99.000 180.825 99.250 181.155 ;
        RECT 99.420 180.865 99.670 181.325 ;
        RECT 96.245 180.385 96.415 180.525 ;
        RECT 95.090 180.345 96.055 180.355 ;
        RECT 94.750 180.175 94.920 180.265 ;
        RECT 95.380 180.185 96.055 180.345 ;
        RECT 92.790 179.985 93.530 180.015 ;
        RECT 92.790 179.685 93.705 179.985 ;
        RECT 93.380 179.510 93.705 179.685 ;
        RECT 92.410 178.955 92.665 179.485 ;
        RECT 92.835 178.775 93.140 179.235 ;
        RECT 93.385 179.155 93.705 179.510 ;
        RECT 93.875 179.725 94.415 180.095 ;
        RECT 94.750 180.005 95.155 180.175 ;
        RECT 93.875 179.325 94.115 179.725 ;
        RECT 94.595 179.555 94.815 179.835 ;
        RECT 94.285 179.385 94.815 179.555 ;
        RECT 94.285 179.155 94.455 179.385 ;
        RECT 94.985 179.225 95.155 180.005 ;
        RECT 95.325 179.395 95.675 180.015 ;
        RECT 95.845 179.395 96.055 180.185 ;
        RECT 96.245 180.215 97.745 180.385 ;
        RECT 96.245 179.525 96.415 180.215 ;
        RECT 98.105 180.045 98.275 180.825 ;
        RECT 99.080 180.695 99.250 180.825 ;
        RECT 96.585 179.875 98.275 180.045 ;
        RECT 98.445 180.265 98.910 180.655 ;
        RECT 99.080 180.525 99.475 180.695 ;
        RECT 96.585 179.695 96.755 179.875 ;
        RECT 93.385 178.985 94.455 179.155 ;
        RECT 94.625 178.775 94.815 179.215 ;
        RECT 94.985 178.945 95.935 179.225 ;
        RECT 96.245 179.135 96.505 179.525 ;
        RECT 96.925 179.455 97.715 179.705 ;
        RECT 96.155 178.965 96.505 179.135 ;
        RECT 96.715 178.775 97.045 179.235 ;
        RECT 97.920 179.165 98.090 179.875 ;
        RECT 98.445 179.675 98.615 180.265 ;
        RECT 98.260 179.455 98.615 179.675 ;
        RECT 98.785 179.455 99.135 180.075 ;
        RECT 99.305 179.165 99.475 180.525 ;
        RECT 99.840 180.355 100.165 181.140 ;
        RECT 99.645 179.305 100.105 180.355 ;
        RECT 97.920 178.995 98.775 179.165 ;
        RECT 98.980 178.995 99.475 179.165 ;
        RECT 99.645 178.775 99.975 179.135 ;
        RECT 100.335 179.035 100.505 181.155 ;
        RECT 100.675 180.825 101.005 181.325 ;
        RECT 101.175 180.655 101.430 181.155 ;
        RECT 100.680 180.485 101.430 180.655 ;
        RECT 100.680 179.495 100.910 180.485 ;
        RECT 101.080 179.665 101.430 180.315 ;
        RECT 101.605 180.160 101.895 181.325 ;
        RECT 102.065 180.185 102.450 181.155 ;
        RECT 102.620 180.865 102.945 181.325 ;
        RECT 103.465 180.695 103.745 181.155 ;
        RECT 102.620 180.475 103.745 180.695 ;
        RECT 102.065 179.515 102.345 180.185 ;
        RECT 102.620 180.015 103.070 180.475 ;
        RECT 103.935 180.305 104.335 181.155 ;
        RECT 104.735 180.865 105.005 181.325 ;
        RECT 105.175 180.695 105.460 181.155 ;
        RECT 102.515 179.685 103.070 180.015 ;
        RECT 103.240 179.745 104.335 180.305 ;
        RECT 102.620 179.575 103.070 179.685 ;
        RECT 100.680 179.325 101.430 179.495 ;
        RECT 100.675 178.775 101.005 179.155 ;
        RECT 101.175 179.035 101.430 179.325 ;
        RECT 101.605 178.775 101.895 179.500 ;
        RECT 102.065 178.945 102.450 179.515 ;
        RECT 102.620 179.405 103.745 179.575 ;
        RECT 102.620 178.775 102.945 179.235 ;
        RECT 103.465 178.945 103.745 179.405 ;
        RECT 103.935 178.945 104.335 179.745 ;
        RECT 104.505 180.475 105.460 180.695 ;
        RECT 104.505 179.575 104.715 180.475 ;
        RECT 104.885 179.745 105.575 180.305 ;
        RECT 105.745 180.185 106.130 181.155 ;
        RECT 106.300 180.865 106.625 181.325 ;
        RECT 107.145 180.695 107.425 181.155 ;
        RECT 106.300 180.475 107.425 180.695 ;
        RECT 104.505 179.405 105.460 179.575 ;
        RECT 104.735 178.775 105.005 179.235 ;
        RECT 105.175 178.945 105.460 179.405 ;
        RECT 105.745 179.515 106.025 180.185 ;
        RECT 106.300 180.015 106.750 180.475 ;
        RECT 107.615 180.305 108.015 181.155 ;
        RECT 108.415 180.865 108.685 181.325 ;
        RECT 108.855 180.695 109.140 181.155 ;
        RECT 106.195 179.685 106.750 180.015 ;
        RECT 106.920 179.745 108.015 180.305 ;
        RECT 106.300 179.575 106.750 179.685 ;
        RECT 105.745 178.945 106.130 179.515 ;
        RECT 106.300 179.405 107.425 179.575 ;
        RECT 106.300 178.775 106.625 179.235 ;
        RECT 107.145 178.945 107.425 179.405 ;
        RECT 107.615 178.945 108.015 179.745 ;
        RECT 108.185 180.475 109.140 180.695 ;
        RECT 108.185 179.575 108.395 180.475 ;
        RECT 108.565 179.745 109.255 180.305 ;
        RECT 109.925 180.185 110.155 181.325 ;
        RECT 110.325 180.175 110.655 181.155 ;
        RECT 110.825 180.185 111.035 181.325 ;
        RECT 109.905 179.765 110.235 180.015 ;
        RECT 108.185 179.405 109.140 179.575 ;
        RECT 108.415 178.775 108.685 179.235 ;
        RECT 108.855 178.945 109.140 179.405 ;
        RECT 109.925 178.775 110.155 179.595 ;
        RECT 110.405 179.575 110.655 180.175 ;
        RECT 111.270 180.135 111.525 181.015 ;
        RECT 111.695 180.185 112.000 181.325 ;
        RECT 112.340 180.945 112.670 181.325 ;
        RECT 112.850 180.775 113.020 181.065 ;
        RECT 113.190 180.865 113.440 181.325 ;
        RECT 112.220 180.605 113.020 180.775 ;
        RECT 113.610 180.815 114.480 181.155 ;
        RECT 110.325 178.945 110.655 179.575 ;
        RECT 110.825 178.775 111.035 179.595 ;
        RECT 111.270 179.485 111.480 180.135 ;
        RECT 112.220 180.015 112.390 180.605 ;
        RECT 113.610 180.435 113.780 180.815 ;
        RECT 114.715 180.695 114.885 181.155 ;
        RECT 115.055 180.865 115.425 181.325 ;
        RECT 115.720 180.725 115.890 181.065 ;
        RECT 116.060 180.895 116.390 181.325 ;
        RECT 116.625 180.725 116.795 181.065 ;
        RECT 112.560 180.265 113.780 180.435 ;
        RECT 113.950 180.355 114.410 180.645 ;
        RECT 114.715 180.525 115.275 180.695 ;
        RECT 115.720 180.555 116.795 180.725 ;
        RECT 116.965 180.825 117.645 181.155 ;
        RECT 117.860 180.825 118.110 181.155 ;
        RECT 118.280 180.865 118.530 181.325 ;
        RECT 115.105 180.385 115.275 180.525 ;
        RECT 113.950 180.345 114.915 180.355 ;
        RECT 113.610 180.175 113.780 180.265 ;
        RECT 114.240 180.185 114.915 180.345 ;
        RECT 111.650 179.985 112.390 180.015 ;
        RECT 111.650 179.685 112.565 179.985 ;
        RECT 112.240 179.510 112.565 179.685 ;
        RECT 111.270 178.955 111.525 179.485 ;
        RECT 111.695 178.775 112.000 179.235 ;
        RECT 112.245 179.155 112.565 179.510 ;
        RECT 112.735 179.725 113.275 180.095 ;
        RECT 113.610 180.005 114.015 180.175 ;
        RECT 112.735 179.325 112.975 179.725 ;
        RECT 113.455 179.555 113.675 179.835 ;
        RECT 113.145 179.385 113.675 179.555 ;
        RECT 113.145 179.155 113.315 179.385 ;
        RECT 113.845 179.225 114.015 180.005 ;
        RECT 114.185 179.395 114.535 180.015 ;
        RECT 114.705 179.395 114.915 180.185 ;
        RECT 115.105 180.215 116.605 180.385 ;
        RECT 115.105 179.525 115.275 180.215 ;
        RECT 116.965 180.045 117.135 180.825 ;
        RECT 117.940 180.695 118.110 180.825 ;
        RECT 115.445 179.875 117.135 180.045 ;
        RECT 117.305 180.265 117.770 180.655 ;
        RECT 117.940 180.525 118.335 180.695 ;
        RECT 115.445 179.695 115.615 179.875 ;
        RECT 112.245 178.985 113.315 179.155 ;
        RECT 113.485 178.775 113.675 179.215 ;
        RECT 113.845 178.945 114.795 179.225 ;
        RECT 115.105 179.135 115.365 179.525 ;
        RECT 115.785 179.455 116.575 179.705 ;
        RECT 115.015 178.965 115.365 179.135 ;
        RECT 115.575 178.775 115.905 179.235 ;
        RECT 116.780 179.165 116.950 179.875 ;
        RECT 117.305 179.675 117.475 180.265 ;
        RECT 117.120 179.455 117.475 179.675 ;
        RECT 117.645 179.455 117.995 180.075 ;
        RECT 118.165 179.165 118.335 180.525 ;
        RECT 118.700 180.355 119.025 181.140 ;
        RECT 118.505 179.305 118.965 180.355 ;
        RECT 116.780 178.995 117.635 179.165 ;
        RECT 117.840 178.995 118.335 179.165 ;
        RECT 118.505 178.775 118.835 179.135 ;
        RECT 119.195 179.035 119.365 181.155 ;
        RECT 119.535 180.825 119.865 181.325 ;
        RECT 120.035 180.655 120.290 181.155 ;
        RECT 119.540 180.485 120.290 180.655 ;
        RECT 119.540 179.495 119.770 180.485 ;
        RECT 119.940 179.665 120.290 180.315 ;
        RECT 120.505 180.185 120.735 181.325 ;
        RECT 120.905 180.175 121.235 181.155 ;
        RECT 121.405 180.185 121.615 181.325 ;
        RECT 121.935 180.395 122.105 181.155 ;
        RECT 122.285 180.565 122.615 181.325 ;
        RECT 121.935 180.225 122.600 180.395 ;
        RECT 122.785 180.250 123.055 181.155 ;
        RECT 120.485 179.765 120.815 180.015 ;
        RECT 119.540 179.325 120.290 179.495 ;
        RECT 119.535 178.775 119.865 179.155 ;
        RECT 120.035 179.035 120.290 179.325 ;
        RECT 120.505 178.775 120.735 179.595 ;
        RECT 120.985 179.575 121.235 180.175 ;
        RECT 122.430 180.080 122.600 180.225 ;
        RECT 121.865 179.675 122.195 180.045 ;
        RECT 122.430 179.750 122.715 180.080 ;
        RECT 120.905 178.945 121.235 179.575 ;
        RECT 121.405 178.775 121.615 179.595 ;
        RECT 122.430 179.495 122.600 179.750 ;
        RECT 121.935 179.325 122.600 179.495 ;
        RECT 122.885 179.450 123.055 180.250 ;
        RECT 123.685 180.235 126.275 181.325 ;
        RECT 126.445 180.235 127.655 181.325 ;
        RECT 123.685 179.715 124.895 180.235 ;
        RECT 125.065 179.545 126.275 180.065 ;
        RECT 126.445 179.695 126.965 180.235 ;
        RECT 121.935 178.945 122.105 179.325 ;
        RECT 122.285 178.775 122.615 179.155 ;
        RECT 122.795 178.945 123.055 179.450 ;
        RECT 123.685 178.775 126.275 179.545 ;
        RECT 127.135 179.525 127.655 180.065 ;
        RECT 126.445 178.775 127.655 179.525 ;
        RECT 14.580 178.605 127.740 178.775 ;
        RECT 14.665 177.855 15.875 178.605 ;
        RECT 14.665 177.315 15.185 177.855 ;
        RECT 16.045 177.835 19.555 178.605 ;
        RECT 19.730 178.060 25.075 178.605 ;
        RECT 15.355 177.145 15.875 177.685 ;
        RECT 14.665 176.055 15.875 177.145 ;
        RECT 16.045 177.145 17.735 177.665 ;
        RECT 17.905 177.315 19.555 177.835 ;
        RECT 16.045 176.055 19.555 177.145 ;
        RECT 21.320 176.490 21.670 177.740 ;
        RECT 23.150 177.230 23.490 178.060 ;
        RECT 25.305 177.785 25.515 178.605 ;
        RECT 25.685 177.805 26.015 178.435 ;
        RECT 25.685 177.205 25.935 177.805 ;
        RECT 26.185 177.785 26.415 178.605 ;
        RECT 26.665 177.785 26.895 178.605 ;
        RECT 27.065 177.805 27.395 178.435 ;
        RECT 26.105 177.365 26.435 177.615 ;
        RECT 26.645 177.365 26.975 177.615 ;
        RECT 27.145 177.205 27.395 177.805 ;
        RECT 27.565 177.785 27.775 178.605 ;
        RECT 28.010 177.895 28.265 178.425 ;
        RECT 28.435 178.145 28.740 178.605 ;
        RECT 28.985 178.225 30.055 178.395 ;
        RECT 19.730 176.055 25.075 176.490 ;
        RECT 25.305 176.055 25.515 177.195 ;
        RECT 25.685 176.225 26.015 177.205 ;
        RECT 26.185 176.055 26.415 177.195 ;
        RECT 26.665 176.055 26.895 177.195 ;
        RECT 27.065 176.225 27.395 177.205 ;
        RECT 28.010 177.245 28.220 177.895 ;
        RECT 28.985 177.870 29.305 178.225 ;
        RECT 28.980 177.695 29.305 177.870 ;
        RECT 28.390 177.395 29.305 177.695 ;
        RECT 29.475 177.655 29.715 178.055 ;
        RECT 29.885 177.995 30.055 178.225 ;
        RECT 30.225 178.165 30.415 178.605 ;
        RECT 30.585 178.155 31.535 178.435 ;
        RECT 31.755 178.245 32.105 178.415 ;
        RECT 29.885 177.825 30.415 177.995 ;
        RECT 28.390 177.365 29.130 177.395 ;
        RECT 27.565 176.055 27.775 177.195 ;
        RECT 28.010 176.365 28.265 177.245 ;
        RECT 28.435 176.055 28.740 177.195 ;
        RECT 28.960 176.775 29.130 177.365 ;
        RECT 29.475 177.285 30.015 177.655 ;
        RECT 30.195 177.545 30.415 177.825 ;
        RECT 30.585 177.375 30.755 178.155 ;
        RECT 30.350 177.205 30.755 177.375 ;
        RECT 30.925 177.365 31.275 177.985 ;
        RECT 30.350 177.115 30.520 177.205 ;
        RECT 31.445 177.195 31.655 177.985 ;
        RECT 29.300 176.945 30.520 177.115 ;
        RECT 30.980 177.035 31.655 177.195 ;
        RECT 28.960 176.605 29.760 176.775 ;
        RECT 29.080 176.055 29.410 176.435 ;
        RECT 29.590 176.315 29.760 176.605 ;
        RECT 30.350 176.565 30.520 176.945 ;
        RECT 30.690 177.025 31.655 177.035 ;
        RECT 31.845 177.855 32.105 178.245 ;
        RECT 32.315 178.145 32.645 178.605 ;
        RECT 33.520 178.215 34.375 178.385 ;
        RECT 34.580 178.215 35.075 178.385 ;
        RECT 35.245 178.245 35.575 178.605 ;
        RECT 31.845 177.165 32.015 177.855 ;
        RECT 32.185 177.505 32.355 177.685 ;
        RECT 32.525 177.675 33.315 177.925 ;
        RECT 33.520 177.505 33.690 178.215 ;
        RECT 33.860 177.705 34.215 177.925 ;
        RECT 32.185 177.335 33.875 177.505 ;
        RECT 30.690 176.735 31.150 177.025 ;
        RECT 31.845 176.995 33.345 177.165 ;
        RECT 31.845 176.855 32.015 176.995 ;
        RECT 31.455 176.685 32.015 176.855 ;
        RECT 29.930 176.055 30.180 176.515 ;
        RECT 30.350 176.225 31.220 176.565 ;
        RECT 31.455 176.225 31.625 176.685 ;
        RECT 32.460 176.655 33.535 176.825 ;
        RECT 31.795 176.055 32.165 176.515 ;
        RECT 32.460 176.315 32.630 176.655 ;
        RECT 32.800 176.055 33.130 176.485 ;
        RECT 33.365 176.315 33.535 176.655 ;
        RECT 33.705 176.555 33.875 177.335 ;
        RECT 34.045 177.115 34.215 177.705 ;
        RECT 34.385 177.305 34.735 177.925 ;
        RECT 34.045 176.725 34.510 177.115 ;
        RECT 34.905 176.855 35.075 178.215 ;
        RECT 35.245 177.025 35.705 178.075 ;
        RECT 34.680 176.685 35.075 176.855 ;
        RECT 34.680 176.555 34.850 176.685 ;
        RECT 33.705 176.225 34.385 176.555 ;
        RECT 34.600 176.225 34.850 176.555 ;
        RECT 35.020 176.055 35.270 176.515 ;
        RECT 35.440 176.240 35.765 177.025 ;
        RECT 35.935 176.225 36.105 178.345 ;
        RECT 36.275 178.225 36.605 178.605 ;
        RECT 36.775 178.055 37.030 178.345 ;
        RECT 36.280 177.885 37.030 178.055 ;
        RECT 36.280 176.895 36.510 177.885 ;
        RECT 37.205 177.880 37.495 178.605 ;
        RECT 37.940 177.795 38.185 178.400 ;
        RECT 38.405 178.070 38.915 178.605 ;
        RECT 36.680 177.065 37.030 177.715 ;
        RECT 37.665 177.625 38.895 177.795 ;
        RECT 36.280 176.725 37.030 176.895 ;
        RECT 36.275 176.055 36.605 176.555 ;
        RECT 36.775 176.225 37.030 176.725 ;
        RECT 37.205 176.055 37.495 177.220 ;
        RECT 37.665 176.815 38.005 177.625 ;
        RECT 38.175 177.060 38.925 177.250 ;
        RECT 37.665 176.405 38.180 176.815 ;
        RECT 38.415 176.055 38.585 176.815 ;
        RECT 38.755 176.395 38.925 177.060 ;
        RECT 39.095 177.075 39.285 178.435 ;
        RECT 39.455 178.265 39.730 178.435 ;
        RECT 39.455 178.095 39.735 178.265 ;
        RECT 39.455 177.275 39.730 178.095 ;
        RECT 39.920 178.070 40.450 178.435 ;
        RECT 40.875 178.205 41.205 178.605 ;
        RECT 40.275 178.035 40.450 178.070 ;
        RECT 39.935 177.075 40.105 177.875 ;
        RECT 39.095 176.905 40.105 177.075 ;
        RECT 40.275 177.865 41.205 178.035 ;
        RECT 41.375 177.865 41.630 178.435 ;
        RECT 40.275 176.735 40.445 177.865 ;
        RECT 41.035 177.695 41.205 177.865 ;
        RECT 39.320 176.565 40.445 176.735 ;
        RECT 40.615 177.365 40.810 177.695 ;
        RECT 41.035 177.365 41.290 177.695 ;
        RECT 40.615 176.395 40.785 177.365 ;
        RECT 41.460 177.195 41.630 177.865 ;
        RECT 42.840 177.975 43.125 178.435 ;
        RECT 43.295 178.145 43.565 178.605 ;
        RECT 42.840 177.805 43.795 177.975 ;
        RECT 38.755 176.225 40.785 176.395 ;
        RECT 40.955 176.055 41.125 177.195 ;
        RECT 41.295 176.225 41.630 177.195 ;
        RECT 42.725 177.075 43.415 177.635 ;
        RECT 43.585 176.905 43.795 177.805 ;
        RECT 42.840 176.685 43.795 176.905 ;
        RECT 43.965 177.635 44.365 178.435 ;
        RECT 44.555 177.975 44.835 178.435 ;
        RECT 45.355 178.145 45.680 178.605 ;
        RECT 44.555 177.805 45.680 177.975 ;
        RECT 45.850 177.865 46.235 178.435 ;
        RECT 45.230 177.695 45.680 177.805 ;
        RECT 43.965 177.075 45.060 177.635 ;
        RECT 45.230 177.365 45.785 177.695 ;
        RECT 42.840 176.225 43.125 176.685 ;
        RECT 43.295 176.055 43.565 176.515 ;
        RECT 43.965 176.225 44.365 177.075 ;
        RECT 45.230 176.905 45.680 177.365 ;
        RECT 45.955 177.195 46.235 177.865 ;
        RECT 46.610 177.825 47.110 178.435 ;
        RECT 46.405 177.365 46.755 177.615 ;
        RECT 46.940 177.195 47.110 177.825 ;
        RECT 47.740 177.955 48.070 178.435 ;
        RECT 48.240 178.145 48.465 178.605 ;
        RECT 48.635 177.955 48.965 178.435 ;
        RECT 47.740 177.785 48.965 177.955 ;
        RECT 49.155 177.805 49.405 178.605 ;
        RECT 49.575 177.805 49.915 178.435 ;
        RECT 50.200 177.975 50.485 178.435 ;
        RECT 50.655 178.145 50.925 178.605 ;
        RECT 50.200 177.805 51.155 177.975 ;
        RECT 47.280 177.415 47.610 177.615 ;
        RECT 47.780 177.415 48.110 177.615 ;
        RECT 48.280 177.415 48.700 177.615 ;
        RECT 48.875 177.445 49.570 177.615 ;
        RECT 48.875 177.195 49.045 177.445 ;
        RECT 49.740 177.195 49.915 177.805 ;
        RECT 44.555 176.685 45.680 176.905 ;
        RECT 44.555 176.225 44.835 176.685 ;
        RECT 45.355 176.055 45.680 176.515 ;
        RECT 45.850 176.225 46.235 177.195 ;
        RECT 46.610 177.025 49.045 177.195 ;
        RECT 46.610 176.225 46.940 177.025 ;
        RECT 47.110 176.055 47.440 176.855 ;
        RECT 47.740 176.225 48.070 177.025 ;
        RECT 48.715 176.055 48.965 176.855 ;
        RECT 49.235 176.055 49.405 177.195 ;
        RECT 49.575 176.225 49.915 177.195 ;
        RECT 50.085 177.075 50.775 177.635 ;
        RECT 50.945 176.905 51.155 177.805 ;
        RECT 50.200 176.685 51.155 176.905 ;
        RECT 51.325 177.635 51.725 178.435 ;
        RECT 51.915 177.975 52.195 178.435 ;
        RECT 52.715 178.145 53.040 178.605 ;
        RECT 51.915 177.805 53.040 177.975 ;
        RECT 53.210 177.865 53.595 178.435 ;
        RECT 52.590 177.695 53.040 177.805 ;
        RECT 51.325 177.075 52.420 177.635 ;
        RECT 52.590 177.365 53.145 177.695 ;
        RECT 50.200 176.225 50.485 176.685 ;
        RECT 50.655 176.055 50.925 176.515 ;
        RECT 51.325 176.225 51.725 177.075 ;
        RECT 52.590 176.905 53.040 177.365 ;
        RECT 53.315 177.195 53.595 177.865 ;
        RECT 51.915 176.685 53.040 176.905 ;
        RECT 51.915 176.225 52.195 176.685 ;
        RECT 52.715 176.055 53.040 176.515 ;
        RECT 53.210 176.225 53.595 177.195 ;
        RECT 53.770 177.895 54.025 178.425 ;
        RECT 54.195 178.145 54.500 178.605 ;
        RECT 54.745 178.225 55.815 178.395 ;
        RECT 53.770 177.245 53.980 177.895 ;
        RECT 54.745 177.870 55.065 178.225 ;
        RECT 54.740 177.695 55.065 177.870 ;
        RECT 54.150 177.395 55.065 177.695 ;
        RECT 55.235 177.655 55.475 178.055 ;
        RECT 55.645 177.995 55.815 178.225 ;
        RECT 55.985 178.165 56.175 178.605 ;
        RECT 56.345 178.155 57.295 178.435 ;
        RECT 57.515 178.245 57.865 178.415 ;
        RECT 55.645 177.825 56.175 177.995 ;
        RECT 54.150 177.365 54.890 177.395 ;
        RECT 53.770 176.365 54.025 177.245 ;
        RECT 54.195 176.055 54.500 177.195 ;
        RECT 54.720 176.775 54.890 177.365 ;
        RECT 55.235 177.285 55.775 177.655 ;
        RECT 55.955 177.545 56.175 177.825 ;
        RECT 56.345 177.375 56.515 178.155 ;
        RECT 56.110 177.205 56.515 177.375 ;
        RECT 56.685 177.365 57.035 177.985 ;
        RECT 56.110 177.115 56.280 177.205 ;
        RECT 57.205 177.195 57.415 177.985 ;
        RECT 55.060 176.945 56.280 177.115 ;
        RECT 56.740 177.035 57.415 177.195 ;
        RECT 54.720 176.605 55.520 176.775 ;
        RECT 54.840 176.055 55.170 176.435 ;
        RECT 55.350 176.315 55.520 176.605 ;
        RECT 56.110 176.565 56.280 176.945 ;
        RECT 56.450 177.025 57.415 177.035 ;
        RECT 57.605 177.855 57.865 178.245 ;
        RECT 58.075 178.145 58.405 178.605 ;
        RECT 59.280 178.215 60.135 178.385 ;
        RECT 60.340 178.215 60.835 178.385 ;
        RECT 61.005 178.245 61.335 178.605 ;
        RECT 57.605 177.165 57.775 177.855 ;
        RECT 57.945 177.505 58.115 177.685 ;
        RECT 58.285 177.675 59.075 177.925 ;
        RECT 59.280 177.505 59.450 178.215 ;
        RECT 59.620 177.705 59.975 177.925 ;
        RECT 57.945 177.335 59.635 177.505 ;
        RECT 56.450 176.735 56.910 177.025 ;
        RECT 57.605 176.995 59.105 177.165 ;
        RECT 57.605 176.855 57.775 176.995 ;
        RECT 57.215 176.685 57.775 176.855 ;
        RECT 55.690 176.055 55.940 176.515 ;
        RECT 56.110 176.225 56.980 176.565 ;
        RECT 57.215 176.225 57.385 176.685 ;
        RECT 58.220 176.655 59.295 176.825 ;
        RECT 57.555 176.055 57.925 176.515 ;
        RECT 58.220 176.315 58.390 176.655 ;
        RECT 58.560 176.055 58.890 176.485 ;
        RECT 59.125 176.315 59.295 176.655 ;
        RECT 59.465 176.555 59.635 177.335 ;
        RECT 59.805 177.115 59.975 177.705 ;
        RECT 60.145 177.305 60.495 177.925 ;
        RECT 59.805 176.725 60.270 177.115 ;
        RECT 60.665 176.855 60.835 178.215 ;
        RECT 61.005 177.025 61.465 178.075 ;
        RECT 60.440 176.685 60.835 176.855 ;
        RECT 60.440 176.555 60.610 176.685 ;
        RECT 59.465 176.225 60.145 176.555 ;
        RECT 60.360 176.225 60.610 176.555 ;
        RECT 60.780 176.055 61.030 176.515 ;
        RECT 61.200 176.240 61.525 177.025 ;
        RECT 61.695 176.225 61.865 178.345 ;
        RECT 62.035 178.225 62.365 178.605 ;
        RECT 62.535 178.055 62.790 178.345 ;
        RECT 62.040 177.885 62.790 178.055 ;
        RECT 62.040 176.895 62.270 177.885 ;
        RECT 62.965 177.880 63.255 178.605 ;
        RECT 63.425 177.930 63.685 178.435 ;
        RECT 63.865 178.225 64.195 178.605 ;
        RECT 64.375 178.055 64.545 178.435 ;
        RECT 62.440 177.065 62.790 177.715 ;
        RECT 62.040 176.725 62.790 176.895 ;
        RECT 62.035 176.055 62.365 176.555 ;
        RECT 62.535 176.225 62.790 176.725 ;
        RECT 62.965 176.055 63.255 177.220 ;
        RECT 63.425 177.130 63.595 177.930 ;
        RECT 63.880 177.885 64.545 178.055 ;
        RECT 63.880 177.630 64.050 177.885 ;
        RECT 64.805 177.835 67.395 178.605 ;
        RECT 63.765 177.300 64.050 177.630 ;
        RECT 64.285 177.335 64.615 177.705 ;
        RECT 63.880 177.155 64.050 177.300 ;
        RECT 63.425 176.225 63.695 177.130 ;
        RECT 63.880 176.985 64.545 177.155 ;
        RECT 63.865 176.055 64.195 176.815 ;
        RECT 64.375 176.225 64.545 176.985 ;
        RECT 64.805 177.145 66.015 177.665 ;
        RECT 66.185 177.315 67.395 177.835 ;
        RECT 67.570 177.765 67.830 178.605 ;
        RECT 68.005 177.860 68.260 178.435 ;
        RECT 68.430 178.225 68.760 178.605 ;
        RECT 68.975 178.055 69.145 178.435 ;
        RECT 68.430 177.885 69.145 178.055 ;
        RECT 69.495 178.055 69.665 178.435 ;
        RECT 69.880 178.225 70.210 178.605 ;
        RECT 69.495 177.885 70.210 178.055 ;
        RECT 64.805 176.055 67.395 177.145 ;
        RECT 67.570 176.055 67.830 177.205 ;
        RECT 68.005 177.130 68.175 177.860 ;
        RECT 68.430 177.695 68.600 177.885 ;
        RECT 68.345 177.365 68.600 177.695 ;
        RECT 68.430 177.155 68.600 177.365 ;
        RECT 68.880 177.335 69.235 177.705 ;
        RECT 69.405 177.335 69.760 177.705 ;
        RECT 70.040 177.695 70.210 177.885 ;
        RECT 70.380 177.860 70.635 178.435 ;
        RECT 70.040 177.365 70.295 177.695 ;
        RECT 70.040 177.155 70.210 177.365 ;
        RECT 68.005 176.225 68.260 177.130 ;
        RECT 68.430 176.985 69.145 177.155 ;
        RECT 68.430 176.055 68.760 176.815 ;
        RECT 68.975 176.225 69.145 176.985 ;
        RECT 69.495 176.985 70.210 177.155 ;
        RECT 70.465 177.130 70.635 177.860 ;
        RECT 70.810 177.765 71.070 178.605 ;
        RECT 71.335 178.055 71.505 178.435 ;
        RECT 71.720 178.225 72.050 178.605 ;
        RECT 71.335 177.885 72.050 178.055 ;
        RECT 71.245 177.335 71.600 177.705 ;
        RECT 71.880 177.695 72.050 177.885 ;
        RECT 72.220 177.860 72.475 178.435 ;
        RECT 71.880 177.365 72.135 177.695 ;
        RECT 69.495 176.225 69.665 176.985 ;
        RECT 69.880 176.055 70.210 176.815 ;
        RECT 70.380 176.225 70.635 177.130 ;
        RECT 70.810 176.055 71.070 177.205 ;
        RECT 71.880 177.155 72.050 177.365 ;
        RECT 71.335 176.985 72.050 177.155 ;
        RECT 72.305 177.130 72.475 177.860 ;
        RECT 72.650 177.765 72.910 178.605 ;
        RECT 73.085 177.845 73.795 178.435 ;
        RECT 74.305 178.075 74.635 178.435 ;
        RECT 74.835 178.245 75.165 178.605 ;
        RECT 75.335 178.075 75.665 178.435 ;
        RECT 74.305 177.865 75.665 178.075 ;
        RECT 71.335 176.225 71.505 176.985 ;
        RECT 71.720 176.055 72.050 176.815 ;
        RECT 72.220 176.225 72.475 177.130 ;
        RECT 72.650 176.055 72.910 177.205 ;
        RECT 73.085 176.875 73.290 177.845 ;
        RECT 76.510 177.825 77.010 178.435 ;
        RECT 73.460 177.075 73.790 177.615 ;
        RECT 73.965 177.365 74.460 177.695 ;
        RECT 74.780 177.365 75.155 177.695 ;
        RECT 75.365 177.365 75.675 177.695 ;
        RECT 76.305 177.365 76.655 177.615 ;
        RECT 73.965 177.075 74.290 177.365 ;
        RECT 74.485 176.875 74.815 177.095 ;
        RECT 73.085 176.645 74.815 176.875 ;
        RECT 73.085 176.225 73.785 176.645 ;
        RECT 73.985 176.055 74.315 176.415 ;
        RECT 74.485 176.245 74.815 176.645 ;
        RECT 74.985 176.440 75.155 177.365 ;
        RECT 76.840 177.195 77.010 177.825 ;
        RECT 77.640 177.955 77.970 178.435 ;
        RECT 78.140 178.145 78.365 178.605 ;
        RECT 78.535 177.955 78.865 178.435 ;
        RECT 77.640 177.785 78.865 177.955 ;
        RECT 79.055 177.805 79.305 178.605 ;
        RECT 79.475 177.805 79.815 178.435 ;
        RECT 77.180 177.415 77.510 177.615 ;
        RECT 77.680 177.415 78.010 177.615 ;
        RECT 78.180 177.415 78.600 177.615 ;
        RECT 78.775 177.445 79.470 177.615 ;
        RECT 78.775 177.195 78.945 177.445 ;
        RECT 79.640 177.245 79.815 177.805 ;
        RECT 79.585 177.195 79.815 177.245 ;
        RECT 75.335 176.055 75.665 177.115 ;
        RECT 76.510 177.025 78.945 177.195 ;
        RECT 76.510 176.225 76.840 177.025 ;
        RECT 77.010 176.055 77.340 176.855 ;
        RECT 77.640 176.225 77.970 177.025 ;
        RECT 78.615 176.055 78.865 176.855 ;
        RECT 79.135 176.055 79.305 177.195 ;
        RECT 79.475 176.225 79.815 177.195 ;
        RECT 79.985 177.805 80.325 178.435 ;
        RECT 80.495 177.805 80.745 178.605 ;
        RECT 80.935 177.955 81.265 178.435 ;
        RECT 81.435 178.145 81.660 178.605 ;
        RECT 81.830 177.955 82.160 178.435 ;
        RECT 79.985 177.755 80.215 177.805 ;
        RECT 80.935 177.785 82.160 177.955 ;
        RECT 82.790 177.825 83.290 178.435 ;
        RECT 83.665 177.855 84.875 178.605 ;
        RECT 79.985 177.195 80.160 177.755 ;
        RECT 80.330 177.445 81.025 177.615 ;
        RECT 80.855 177.195 81.025 177.445 ;
        RECT 81.200 177.415 81.620 177.615 ;
        RECT 81.790 177.415 82.120 177.615 ;
        RECT 82.290 177.415 82.620 177.615 ;
        RECT 82.790 177.195 82.960 177.825 ;
        RECT 83.145 177.365 83.495 177.615 ;
        RECT 79.985 176.225 80.325 177.195 ;
        RECT 80.495 176.055 80.665 177.195 ;
        RECT 80.855 177.025 83.290 177.195 ;
        RECT 80.935 176.055 81.185 176.855 ;
        RECT 81.830 176.225 82.160 177.025 ;
        RECT 82.460 176.055 82.790 176.855 ;
        RECT 82.960 176.225 83.290 177.025 ;
        RECT 83.665 177.145 84.185 177.685 ;
        RECT 84.355 177.315 84.875 177.855 ;
        RECT 85.160 177.975 85.445 178.435 ;
        RECT 85.615 178.145 85.885 178.605 ;
        RECT 85.160 177.805 86.115 177.975 ;
        RECT 83.665 176.055 84.875 177.145 ;
        RECT 85.045 177.075 85.735 177.635 ;
        RECT 85.905 176.905 86.115 177.805 ;
        RECT 85.160 176.685 86.115 176.905 ;
        RECT 86.285 177.635 86.685 178.435 ;
        RECT 86.875 177.975 87.155 178.435 ;
        RECT 87.675 178.145 88.000 178.605 ;
        RECT 86.875 177.805 88.000 177.975 ;
        RECT 88.170 177.865 88.555 178.435 ;
        RECT 88.725 177.880 89.015 178.605 ;
        RECT 87.550 177.695 88.000 177.805 ;
        RECT 86.285 177.075 87.380 177.635 ;
        RECT 87.550 177.365 88.105 177.695 ;
        RECT 85.160 176.225 85.445 176.685 ;
        RECT 85.615 176.055 85.885 176.515 ;
        RECT 86.285 176.225 86.685 177.075 ;
        RECT 87.550 176.905 88.000 177.365 ;
        RECT 88.275 177.195 88.555 177.865 ;
        RECT 89.185 177.835 92.695 178.605 ;
        RECT 92.870 178.060 98.215 178.605 ;
        RECT 86.875 176.685 88.000 176.905 ;
        RECT 86.875 176.225 87.155 176.685 ;
        RECT 87.675 176.055 88.000 176.515 ;
        RECT 88.170 176.225 88.555 177.195 ;
        RECT 88.725 176.055 89.015 177.220 ;
        RECT 89.185 177.145 90.875 177.665 ;
        RECT 91.045 177.315 92.695 177.835 ;
        RECT 89.185 176.055 92.695 177.145 ;
        RECT 94.460 176.490 94.810 177.740 ;
        RECT 96.290 177.230 96.630 178.060 ;
        RECT 98.590 177.825 99.090 178.435 ;
        RECT 98.385 177.365 98.735 177.615 ;
        RECT 98.920 177.195 99.090 177.825 ;
        RECT 99.720 177.955 100.050 178.435 ;
        RECT 100.220 178.145 100.445 178.605 ;
        RECT 100.615 177.955 100.945 178.435 ;
        RECT 99.720 177.785 100.945 177.955 ;
        RECT 101.135 177.805 101.385 178.605 ;
        RECT 101.555 177.805 101.895 178.435 ;
        RECT 99.260 177.415 99.590 177.615 ;
        RECT 99.760 177.415 100.090 177.615 ;
        RECT 100.260 177.415 100.680 177.615 ;
        RECT 100.855 177.445 101.550 177.615 ;
        RECT 100.855 177.195 101.025 177.445 ;
        RECT 101.720 177.195 101.895 177.805 ;
        RECT 98.590 177.025 101.025 177.195 ;
        RECT 92.870 176.055 98.215 176.490 ;
        RECT 98.590 176.225 98.920 177.025 ;
        RECT 99.090 176.055 99.420 176.855 ;
        RECT 99.720 176.225 100.050 177.025 ;
        RECT 100.695 176.055 100.945 176.855 ;
        RECT 101.215 176.055 101.385 177.195 ;
        RECT 101.555 176.225 101.895 177.195 ;
        RECT 102.065 177.930 102.325 178.435 ;
        RECT 102.505 178.225 102.835 178.605 ;
        RECT 103.015 178.055 103.185 178.435 ;
        RECT 102.065 177.130 102.235 177.930 ;
        RECT 102.520 177.885 103.185 178.055 ;
        RECT 102.520 177.630 102.690 177.885 ;
        RECT 103.445 177.855 104.655 178.605 ;
        RECT 102.405 177.300 102.690 177.630 ;
        RECT 102.925 177.335 103.255 177.705 ;
        RECT 102.520 177.155 102.690 177.300 ;
        RECT 102.065 176.225 102.335 177.130 ;
        RECT 102.520 176.985 103.185 177.155 ;
        RECT 102.505 176.055 102.835 176.815 ;
        RECT 103.015 176.225 103.185 176.985 ;
        RECT 103.445 177.145 103.965 177.685 ;
        RECT 104.135 177.315 104.655 177.855 ;
        RECT 104.825 177.805 105.165 178.435 ;
        RECT 105.335 177.805 105.585 178.605 ;
        RECT 105.775 177.955 106.105 178.435 ;
        RECT 106.275 178.145 106.500 178.605 ;
        RECT 106.670 177.955 107.000 178.435 ;
        RECT 104.825 177.195 105.000 177.805 ;
        RECT 105.775 177.785 107.000 177.955 ;
        RECT 107.630 177.825 108.130 178.435 ;
        RECT 108.505 177.835 110.175 178.605 ;
        RECT 105.170 177.445 105.865 177.615 ;
        RECT 105.695 177.195 105.865 177.445 ;
        RECT 106.040 177.415 106.460 177.615 ;
        RECT 106.630 177.415 106.960 177.615 ;
        RECT 107.130 177.415 107.460 177.615 ;
        RECT 107.630 177.195 107.800 177.825 ;
        RECT 107.985 177.365 108.335 177.615 ;
        RECT 103.445 176.055 104.655 177.145 ;
        RECT 104.825 176.225 105.165 177.195 ;
        RECT 105.335 176.055 105.505 177.195 ;
        RECT 105.695 177.025 108.130 177.195 ;
        RECT 105.775 176.055 106.025 176.855 ;
        RECT 106.670 176.225 107.000 177.025 ;
        RECT 107.300 176.055 107.630 176.855 ;
        RECT 107.800 176.225 108.130 177.025 ;
        RECT 108.505 177.145 109.255 177.665 ;
        RECT 109.425 177.315 110.175 177.835 ;
        RECT 110.620 177.795 110.865 178.400 ;
        RECT 111.085 178.070 111.595 178.605 ;
        RECT 110.345 177.625 111.575 177.795 ;
        RECT 108.505 176.055 110.175 177.145 ;
        RECT 110.345 176.815 110.685 177.625 ;
        RECT 110.855 177.060 111.605 177.250 ;
        RECT 110.345 176.405 110.860 176.815 ;
        RECT 111.095 176.055 111.265 176.815 ;
        RECT 111.435 176.395 111.605 177.060 ;
        RECT 111.775 177.075 111.965 178.435 ;
        RECT 112.135 178.265 112.410 178.435 ;
        RECT 112.135 178.095 112.415 178.265 ;
        RECT 112.135 177.275 112.410 178.095 ;
        RECT 112.600 178.070 113.130 178.435 ;
        RECT 113.555 178.205 113.885 178.605 ;
        RECT 112.955 178.035 113.130 178.070 ;
        RECT 112.615 177.075 112.785 177.875 ;
        RECT 111.775 176.905 112.785 177.075 ;
        RECT 112.955 177.865 113.885 178.035 ;
        RECT 114.055 177.865 114.310 178.435 ;
        RECT 114.485 177.880 114.775 178.605 ;
        RECT 112.955 176.735 113.125 177.865 ;
        RECT 113.715 177.695 113.885 177.865 ;
        RECT 112.000 176.565 113.125 176.735 ;
        RECT 113.295 177.365 113.490 177.695 ;
        RECT 113.715 177.365 113.970 177.695 ;
        RECT 113.295 176.395 113.465 177.365 ;
        RECT 114.140 177.195 114.310 177.865 ;
        RECT 114.945 177.835 116.615 178.605 ;
        RECT 116.875 178.055 117.045 178.435 ;
        RECT 117.225 178.225 117.555 178.605 ;
        RECT 116.875 177.885 117.540 178.055 ;
        RECT 117.735 177.930 117.995 178.435 ;
        RECT 111.435 176.225 113.465 176.395 ;
        RECT 113.635 176.055 113.805 177.195 ;
        RECT 113.975 176.225 114.310 177.195 ;
        RECT 114.485 176.055 114.775 177.220 ;
        RECT 114.945 177.145 115.695 177.665 ;
        RECT 115.865 177.315 116.615 177.835 ;
        RECT 116.805 177.335 117.135 177.705 ;
        RECT 117.370 177.630 117.540 177.885 ;
        RECT 117.370 177.300 117.655 177.630 ;
        RECT 117.370 177.155 117.540 177.300 ;
        RECT 114.945 176.055 116.615 177.145 ;
        RECT 116.875 176.985 117.540 177.155 ;
        RECT 117.825 177.130 117.995 177.930 ;
        RECT 118.165 177.835 120.755 178.605 ;
        RECT 120.930 178.060 126.275 178.605 ;
        RECT 116.875 176.225 117.045 176.985 ;
        RECT 117.225 176.055 117.555 176.815 ;
        RECT 117.725 176.225 117.995 177.130 ;
        RECT 118.165 177.145 119.375 177.665 ;
        RECT 119.545 177.315 120.755 177.835 ;
        RECT 118.165 176.055 120.755 177.145 ;
        RECT 122.520 176.490 122.870 177.740 ;
        RECT 124.350 177.230 124.690 178.060 ;
        RECT 126.445 177.855 127.655 178.605 ;
        RECT 126.445 177.145 126.965 177.685 ;
        RECT 127.135 177.315 127.655 177.855 ;
        RECT 120.930 176.055 126.275 176.490 ;
        RECT 126.445 176.055 127.655 177.145 ;
        RECT 14.580 175.885 127.740 176.055 ;
        RECT 14.665 174.795 15.875 175.885 ;
        RECT 14.665 174.085 15.185 174.625 ;
        RECT 15.355 174.255 15.875 174.795 ;
        RECT 16.045 174.795 18.635 175.885 ;
        RECT 18.810 175.450 24.155 175.885 ;
        RECT 16.045 174.275 17.255 174.795 ;
        RECT 17.425 174.105 18.635 174.625 ;
        RECT 20.400 174.200 20.750 175.450 ;
        RECT 24.325 174.720 24.615 175.885 ;
        RECT 25.705 174.810 25.975 175.715 ;
        RECT 26.145 175.125 26.475 175.885 ;
        RECT 26.655 174.955 26.825 175.715 ;
        RECT 27.200 175.255 27.485 175.715 ;
        RECT 27.655 175.425 27.925 175.885 ;
        RECT 27.200 175.035 28.155 175.255 ;
        RECT 14.665 173.335 15.875 174.085 ;
        RECT 16.045 173.335 18.635 174.105 ;
        RECT 22.230 173.880 22.570 174.710 ;
        RECT 18.810 173.335 24.155 173.880 ;
        RECT 24.325 173.335 24.615 174.060 ;
        RECT 25.705 174.010 25.875 174.810 ;
        RECT 26.160 174.785 26.825 174.955 ;
        RECT 26.160 174.640 26.330 174.785 ;
        RECT 26.045 174.310 26.330 174.640 ;
        RECT 26.160 174.055 26.330 174.310 ;
        RECT 26.565 174.235 26.895 174.605 ;
        RECT 27.085 174.305 27.775 174.865 ;
        RECT 27.945 174.135 28.155 175.035 ;
        RECT 25.705 173.505 25.965 174.010 ;
        RECT 26.160 173.885 26.825 174.055 ;
        RECT 26.145 173.335 26.475 173.715 ;
        RECT 26.655 173.505 26.825 173.885 ;
        RECT 27.200 173.965 28.155 174.135 ;
        RECT 28.325 174.865 28.725 175.715 ;
        RECT 28.915 175.255 29.195 175.715 ;
        RECT 29.715 175.425 30.040 175.885 ;
        RECT 28.915 175.035 30.040 175.255 ;
        RECT 28.325 174.305 29.420 174.865 ;
        RECT 29.590 174.575 30.040 175.035 ;
        RECT 30.210 174.745 30.595 175.715 ;
        RECT 27.200 173.505 27.485 173.965 ;
        RECT 27.655 173.335 27.925 173.795 ;
        RECT 28.325 173.505 28.725 174.305 ;
        RECT 29.590 174.245 30.145 174.575 ;
        RECT 29.590 174.135 30.040 174.245 ;
        RECT 28.915 173.965 30.040 174.135 ;
        RECT 30.315 174.075 30.595 174.745 ;
        RECT 28.915 173.505 29.195 173.965 ;
        RECT 29.715 173.335 30.040 173.795 ;
        RECT 30.210 173.505 30.595 174.075 ;
        RECT 30.770 174.745 31.105 175.715 ;
        RECT 31.275 174.745 31.445 175.885 ;
        RECT 31.615 175.545 33.645 175.715 ;
        RECT 30.770 174.075 30.940 174.745 ;
        RECT 31.615 174.575 31.785 175.545 ;
        RECT 31.110 174.245 31.365 174.575 ;
        RECT 31.590 174.245 31.785 174.575 ;
        RECT 31.955 175.205 33.080 175.375 ;
        RECT 31.195 174.075 31.365 174.245 ;
        RECT 31.955 174.075 32.125 175.205 ;
        RECT 30.770 173.505 31.025 174.075 ;
        RECT 31.195 173.905 32.125 174.075 ;
        RECT 32.295 174.865 33.305 175.035 ;
        RECT 32.295 174.065 32.465 174.865 ;
        RECT 32.670 174.525 32.945 174.665 ;
        RECT 32.665 174.355 32.945 174.525 ;
        RECT 31.950 173.870 32.125 173.905 ;
        RECT 31.195 173.335 31.525 173.735 ;
        RECT 31.950 173.505 32.480 173.870 ;
        RECT 32.670 173.505 32.945 174.355 ;
        RECT 33.115 173.505 33.305 174.865 ;
        RECT 33.475 174.880 33.645 175.545 ;
        RECT 33.815 175.125 33.985 175.885 ;
        RECT 34.220 175.125 34.735 175.535 ;
        RECT 33.475 174.690 34.225 174.880 ;
        RECT 34.395 174.315 34.735 175.125 ;
        RECT 35.570 174.915 35.900 175.715 ;
        RECT 36.070 175.085 36.400 175.885 ;
        RECT 36.700 174.915 37.030 175.715 ;
        RECT 37.675 175.085 37.925 175.885 ;
        RECT 35.570 174.745 38.005 174.915 ;
        RECT 38.195 174.745 38.365 175.885 ;
        RECT 38.535 174.745 38.875 175.715 ;
        RECT 35.365 174.325 35.715 174.575 ;
        RECT 33.505 174.145 34.735 174.315 ;
        RECT 33.485 173.335 33.995 173.870 ;
        RECT 34.215 173.540 34.460 174.145 ;
        RECT 35.900 174.115 36.070 174.745 ;
        RECT 36.240 174.325 36.570 174.525 ;
        RECT 36.740 174.325 37.070 174.525 ;
        RECT 37.240 174.325 37.660 174.525 ;
        RECT 37.835 174.495 38.005 174.745 ;
        RECT 37.835 174.325 38.530 174.495 ;
        RECT 38.700 174.185 38.875 174.745 ;
        RECT 35.570 173.505 36.070 174.115 ;
        RECT 36.700 173.985 37.925 174.155 ;
        RECT 38.645 174.135 38.875 174.185 ;
        RECT 36.700 173.505 37.030 173.985 ;
        RECT 37.200 173.335 37.425 173.795 ;
        RECT 37.595 173.505 37.925 173.985 ;
        RECT 38.115 173.335 38.365 174.135 ;
        RECT 38.535 173.505 38.875 174.135 ;
        RECT 39.045 174.745 39.385 175.715 ;
        RECT 39.555 174.745 39.725 175.885 ;
        RECT 39.995 175.085 40.245 175.885 ;
        RECT 40.890 174.915 41.220 175.715 ;
        RECT 41.520 175.085 41.850 175.885 ;
        RECT 42.020 174.915 42.350 175.715 ;
        RECT 39.915 174.745 42.350 174.915 ;
        RECT 42.930 174.915 43.260 175.715 ;
        RECT 43.430 175.085 43.760 175.885 ;
        RECT 44.060 174.915 44.390 175.715 ;
        RECT 45.035 175.085 45.285 175.885 ;
        RECT 42.930 174.745 45.365 174.915 ;
        RECT 45.555 174.745 45.725 175.885 ;
        RECT 45.895 174.745 46.235 175.715 ;
        RECT 46.520 175.255 46.805 175.715 ;
        RECT 46.975 175.425 47.245 175.885 ;
        RECT 46.520 175.035 47.475 175.255 ;
        RECT 39.045 174.135 39.220 174.745 ;
        RECT 39.915 174.495 40.085 174.745 ;
        RECT 39.390 174.325 40.085 174.495 ;
        RECT 40.260 174.325 40.680 174.525 ;
        RECT 40.850 174.325 41.180 174.525 ;
        RECT 41.350 174.325 41.680 174.525 ;
        RECT 39.045 173.505 39.385 174.135 ;
        RECT 39.555 173.335 39.805 174.135 ;
        RECT 39.995 173.985 41.220 174.155 ;
        RECT 39.995 173.505 40.325 173.985 ;
        RECT 40.495 173.335 40.720 173.795 ;
        RECT 40.890 173.505 41.220 173.985 ;
        RECT 41.850 174.115 42.020 174.745 ;
        RECT 42.205 174.325 42.555 174.575 ;
        RECT 42.725 174.325 43.075 174.575 ;
        RECT 43.260 174.115 43.430 174.745 ;
        RECT 43.600 174.325 43.930 174.525 ;
        RECT 44.100 174.325 44.430 174.525 ;
        RECT 44.600 174.325 45.020 174.525 ;
        RECT 45.195 174.495 45.365 174.745 ;
        RECT 45.195 174.325 45.890 174.495 ;
        RECT 46.060 174.185 46.235 174.745 ;
        RECT 46.405 174.305 47.095 174.865 ;
        RECT 41.850 173.505 42.350 174.115 ;
        RECT 42.930 173.505 43.430 174.115 ;
        RECT 44.060 173.985 45.285 174.155 ;
        RECT 46.005 174.135 46.235 174.185 ;
        RECT 47.265 174.135 47.475 175.035 ;
        RECT 44.060 173.505 44.390 173.985 ;
        RECT 44.560 173.335 44.785 173.795 ;
        RECT 44.955 173.505 45.285 173.985 ;
        RECT 45.475 173.335 45.725 174.135 ;
        RECT 45.895 173.505 46.235 174.135 ;
        RECT 46.520 173.965 47.475 174.135 ;
        RECT 47.645 174.865 48.045 175.715 ;
        RECT 48.235 175.255 48.515 175.715 ;
        RECT 49.035 175.425 49.360 175.885 ;
        RECT 48.235 175.035 49.360 175.255 ;
        RECT 47.645 174.305 48.740 174.865 ;
        RECT 48.910 174.575 49.360 175.035 ;
        RECT 49.530 174.745 49.915 175.715 ;
        RECT 46.520 173.505 46.805 173.965 ;
        RECT 46.975 173.335 47.245 173.795 ;
        RECT 47.645 173.505 48.045 174.305 ;
        RECT 48.910 174.245 49.465 174.575 ;
        RECT 48.910 174.135 49.360 174.245 ;
        RECT 48.235 173.965 49.360 174.135 ;
        RECT 49.635 174.075 49.915 174.745 ;
        RECT 50.085 174.720 50.375 175.885 ;
        RECT 50.545 174.795 53.135 175.885 ;
        RECT 53.305 175.125 53.820 175.535 ;
        RECT 54.055 175.125 54.225 175.885 ;
        RECT 54.395 175.545 56.425 175.715 ;
        RECT 50.545 174.275 51.755 174.795 ;
        RECT 51.925 174.105 53.135 174.625 ;
        RECT 53.305 174.315 53.645 175.125 ;
        RECT 54.395 174.880 54.565 175.545 ;
        RECT 54.960 175.205 56.085 175.375 ;
        RECT 53.815 174.690 54.565 174.880 ;
        RECT 54.735 174.865 55.745 175.035 ;
        RECT 53.305 174.145 54.535 174.315 ;
        RECT 48.235 173.505 48.515 173.965 ;
        RECT 49.035 173.335 49.360 173.795 ;
        RECT 49.530 173.505 49.915 174.075 ;
        RECT 50.085 173.335 50.375 174.060 ;
        RECT 50.545 173.335 53.135 174.105 ;
        RECT 53.580 173.540 53.825 174.145 ;
        RECT 54.045 173.335 54.555 173.870 ;
        RECT 54.735 173.505 54.925 174.865 ;
        RECT 55.095 174.525 55.370 174.665 ;
        RECT 55.095 174.355 55.375 174.525 ;
        RECT 55.095 173.505 55.370 174.355 ;
        RECT 55.575 174.065 55.745 174.865 ;
        RECT 55.915 174.075 56.085 175.205 ;
        RECT 56.255 174.575 56.425 175.545 ;
        RECT 56.595 174.745 56.765 175.885 ;
        RECT 56.935 174.745 57.270 175.715 ;
        RECT 56.255 174.245 56.450 174.575 ;
        RECT 56.675 174.245 56.930 174.575 ;
        RECT 56.675 174.075 56.845 174.245 ;
        RECT 57.100 174.075 57.270 174.745 ;
        RECT 55.915 173.905 56.845 174.075 ;
        RECT 55.915 173.870 56.090 173.905 ;
        RECT 55.560 173.505 56.090 173.870 ;
        RECT 56.515 173.335 56.845 173.735 ;
        RECT 57.015 173.505 57.270 174.075 ;
        RECT 57.450 174.695 57.705 175.575 ;
        RECT 57.875 174.745 58.180 175.885 ;
        RECT 58.520 175.505 58.850 175.885 ;
        RECT 59.030 175.335 59.200 175.625 ;
        RECT 59.370 175.425 59.620 175.885 ;
        RECT 58.400 175.165 59.200 175.335 ;
        RECT 59.790 175.375 60.660 175.715 ;
        RECT 57.450 174.045 57.660 174.695 ;
        RECT 58.400 174.575 58.570 175.165 ;
        RECT 59.790 174.995 59.960 175.375 ;
        RECT 60.895 175.255 61.065 175.715 ;
        RECT 61.235 175.425 61.605 175.885 ;
        RECT 61.900 175.285 62.070 175.625 ;
        RECT 62.240 175.455 62.570 175.885 ;
        RECT 62.805 175.285 62.975 175.625 ;
        RECT 58.740 174.825 59.960 174.995 ;
        RECT 60.130 174.915 60.590 175.205 ;
        RECT 60.895 175.085 61.455 175.255 ;
        RECT 61.900 175.115 62.975 175.285 ;
        RECT 63.145 175.385 63.825 175.715 ;
        RECT 64.040 175.385 64.290 175.715 ;
        RECT 64.460 175.425 64.710 175.885 ;
        RECT 61.285 174.945 61.455 175.085 ;
        RECT 60.130 174.905 61.095 174.915 ;
        RECT 59.790 174.735 59.960 174.825 ;
        RECT 60.420 174.745 61.095 174.905 ;
        RECT 57.830 174.545 58.570 174.575 ;
        RECT 57.830 174.245 58.745 174.545 ;
        RECT 58.420 174.070 58.745 174.245 ;
        RECT 57.450 173.515 57.705 174.045 ;
        RECT 57.875 173.335 58.180 173.795 ;
        RECT 58.425 173.715 58.745 174.070 ;
        RECT 58.915 174.285 59.455 174.655 ;
        RECT 59.790 174.565 60.195 174.735 ;
        RECT 58.915 173.885 59.155 174.285 ;
        RECT 59.635 174.115 59.855 174.395 ;
        RECT 59.325 173.945 59.855 174.115 ;
        RECT 59.325 173.715 59.495 173.945 ;
        RECT 60.025 173.785 60.195 174.565 ;
        RECT 60.365 173.955 60.715 174.575 ;
        RECT 60.885 173.955 61.095 174.745 ;
        RECT 61.285 174.775 62.785 174.945 ;
        RECT 61.285 174.085 61.455 174.775 ;
        RECT 63.145 174.605 63.315 175.385 ;
        RECT 64.120 175.255 64.290 175.385 ;
        RECT 61.625 174.435 63.315 174.605 ;
        RECT 63.485 174.825 63.950 175.215 ;
        RECT 64.120 175.085 64.515 175.255 ;
        RECT 61.625 174.255 61.795 174.435 ;
        RECT 58.425 173.545 59.495 173.715 ;
        RECT 59.665 173.335 59.855 173.775 ;
        RECT 60.025 173.505 60.975 173.785 ;
        RECT 61.285 173.695 61.545 174.085 ;
        RECT 61.965 174.015 62.755 174.265 ;
        RECT 61.195 173.525 61.545 173.695 ;
        RECT 61.755 173.335 62.085 173.795 ;
        RECT 62.960 173.725 63.130 174.435 ;
        RECT 63.485 174.235 63.655 174.825 ;
        RECT 63.300 174.015 63.655 174.235 ;
        RECT 63.825 174.015 64.175 174.635 ;
        RECT 64.345 173.725 64.515 175.085 ;
        RECT 64.880 174.915 65.205 175.700 ;
        RECT 64.685 173.865 65.145 174.915 ;
        RECT 62.960 173.555 63.815 173.725 ;
        RECT 64.020 173.555 64.515 173.725 ;
        RECT 64.685 173.335 65.015 173.695 ;
        RECT 65.375 173.595 65.545 175.715 ;
        RECT 65.715 175.385 66.045 175.885 ;
        RECT 66.215 175.215 66.470 175.715 ;
        RECT 65.720 175.045 66.470 175.215 ;
        RECT 65.720 174.055 65.950 175.045 ;
        RECT 66.120 174.225 66.470 174.875 ;
        RECT 66.645 174.795 68.315 175.885 ;
        RECT 68.495 174.905 68.825 175.715 ;
        RECT 68.995 175.085 69.235 175.885 ;
        RECT 66.645 174.275 67.395 174.795 ;
        RECT 68.495 174.735 69.210 174.905 ;
        RECT 67.565 174.105 68.315 174.625 ;
        RECT 68.490 174.325 68.870 174.565 ;
        RECT 69.040 174.495 69.210 174.735 ;
        RECT 69.415 174.865 69.585 175.715 ;
        RECT 69.755 175.085 70.085 175.885 ;
        RECT 70.255 174.865 70.425 175.715 ;
        RECT 69.415 174.695 70.425 174.865 ;
        RECT 70.595 174.735 70.925 175.885 ;
        RECT 71.250 174.735 71.510 175.885 ;
        RECT 71.685 174.810 71.940 175.715 ;
        RECT 72.110 175.125 72.440 175.885 ;
        RECT 72.655 174.955 72.825 175.715 ;
        RECT 69.040 174.325 69.540 174.495 ;
        RECT 69.040 174.155 69.210 174.325 ;
        RECT 69.930 174.155 70.425 174.695 ;
        RECT 65.720 173.885 66.470 174.055 ;
        RECT 65.715 173.335 66.045 173.715 ;
        RECT 66.215 173.595 66.470 173.885 ;
        RECT 66.645 173.335 68.315 174.105 ;
        RECT 68.575 173.985 69.210 174.155 ;
        RECT 69.415 173.985 70.425 174.155 ;
        RECT 68.575 173.505 68.745 173.985 ;
        RECT 68.925 173.335 69.165 173.815 ;
        RECT 69.415 173.505 69.585 173.985 ;
        RECT 69.755 173.335 70.085 173.815 ;
        RECT 70.255 173.505 70.425 173.985 ;
        RECT 70.595 173.335 70.925 174.135 ;
        RECT 71.250 173.335 71.510 174.175 ;
        RECT 71.685 174.080 71.855 174.810 ;
        RECT 72.110 174.785 72.825 174.955 ;
        RECT 73.085 174.795 75.675 175.885 ;
        RECT 72.110 174.575 72.280 174.785 ;
        RECT 72.025 174.245 72.280 174.575 ;
        RECT 71.685 173.505 71.940 174.080 ;
        RECT 72.110 174.055 72.280 174.245 ;
        RECT 72.560 174.235 72.915 174.605 ;
        RECT 73.085 174.275 74.295 174.795 ;
        RECT 75.845 174.720 76.135 175.885 ;
        RECT 77.225 174.795 80.735 175.885 ;
        RECT 74.465 174.105 75.675 174.625 ;
        RECT 77.225 174.275 78.915 174.795 ;
        RECT 80.905 174.745 81.245 175.715 ;
        RECT 81.415 174.745 81.585 175.885 ;
        RECT 81.855 175.085 82.105 175.885 ;
        RECT 82.750 174.915 83.080 175.715 ;
        RECT 83.380 175.085 83.710 175.885 ;
        RECT 83.880 174.915 84.210 175.715 ;
        RECT 85.050 175.450 90.395 175.885 ;
        RECT 90.570 175.450 95.915 175.885 ;
        RECT 96.090 175.450 101.435 175.885 ;
        RECT 81.775 174.745 84.210 174.915 ;
        RECT 79.085 174.105 80.735 174.625 ;
        RECT 72.110 173.885 72.825 174.055 ;
        RECT 72.110 173.335 72.440 173.715 ;
        RECT 72.655 173.505 72.825 173.885 ;
        RECT 73.085 173.335 75.675 174.105 ;
        RECT 75.845 173.335 76.135 174.060 ;
        RECT 77.225 173.335 80.735 174.105 ;
        RECT 80.905 174.185 81.080 174.745 ;
        RECT 81.775 174.495 81.945 174.745 ;
        RECT 81.250 174.325 81.945 174.495 ;
        RECT 82.120 174.325 82.540 174.525 ;
        RECT 82.710 174.325 83.040 174.525 ;
        RECT 83.210 174.325 83.540 174.525 ;
        RECT 80.905 174.135 81.135 174.185 ;
        RECT 80.905 173.505 81.245 174.135 ;
        RECT 81.415 173.335 81.665 174.135 ;
        RECT 81.855 173.985 83.080 174.155 ;
        RECT 81.855 173.505 82.185 173.985 ;
        RECT 82.355 173.335 82.580 173.795 ;
        RECT 82.750 173.505 83.080 173.985 ;
        RECT 83.710 174.115 83.880 174.745 ;
        RECT 84.065 174.325 84.415 174.575 ;
        RECT 86.640 174.200 86.990 175.450 ;
        RECT 83.710 173.505 84.210 174.115 ;
        RECT 88.470 173.880 88.810 174.710 ;
        RECT 92.160 174.200 92.510 175.450 ;
        RECT 93.990 173.880 94.330 174.710 ;
        RECT 97.680 174.200 98.030 175.450 ;
        RECT 101.605 174.720 101.895 175.885 ;
        RECT 102.065 174.795 103.735 175.885 ;
        RECT 104.110 174.915 104.440 175.715 ;
        RECT 104.610 175.085 104.940 175.885 ;
        RECT 105.240 174.915 105.570 175.715 ;
        RECT 106.215 175.085 106.465 175.885 ;
        RECT 99.510 173.880 99.850 174.710 ;
        RECT 102.065 174.275 102.815 174.795 ;
        RECT 104.110 174.745 106.545 174.915 ;
        RECT 106.735 174.745 106.905 175.885 ;
        RECT 107.075 174.745 107.415 175.715 ;
        RECT 102.985 174.105 103.735 174.625 ;
        RECT 103.905 174.325 104.255 174.575 ;
        RECT 104.440 174.115 104.610 174.745 ;
        RECT 104.780 174.325 105.110 174.525 ;
        RECT 105.280 174.325 105.610 174.525 ;
        RECT 105.780 174.325 106.200 174.525 ;
        RECT 106.375 174.495 106.545 174.745 ;
        RECT 106.375 174.325 107.070 174.495 ;
        RECT 85.050 173.335 90.395 173.880 ;
        RECT 90.570 173.335 95.915 173.880 ;
        RECT 96.090 173.335 101.435 173.880 ;
        RECT 101.605 173.335 101.895 174.060 ;
        RECT 102.065 173.335 103.735 174.105 ;
        RECT 104.110 173.505 104.610 174.115 ;
        RECT 105.240 173.985 106.465 174.155 ;
        RECT 107.240 174.135 107.415 174.745 ;
        RECT 105.240 173.505 105.570 173.985 ;
        RECT 105.740 173.335 105.965 173.795 ;
        RECT 106.135 173.505 106.465 173.985 ;
        RECT 106.655 173.335 106.905 174.135 ;
        RECT 107.075 173.505 107.415 174.135 ;
        RECT 107.585 174.745 107.925 175.715 ;
        RECT 108.095 174.745 108.265 175.885 ;
        RECT 108.535 175.085 108.785 175.885 ;
        RECT 109.430 174.915 109.760 175.715 ;
        RECT 110.060 175.085 110.390 175.885 ;
        RECT 110.560 174.915 110.890 175.715 ;
        RECT 108.455 174.745 110.890 174.915 ;
        RECT 111.265 174.795 112.475 175.885 ;
        RECT 112.650 175.450 117.995 175.885 ;
        RECT 107.585 174.185 107.760 174.745 ;
        RECT 108.455 174.495 108.625 174.745 ;
        RECT 107.930 174.325 108.625 174.495 ;
        RECT 108.800 174.325 109.220 174.525 ;
        RECT 109.390 174.325 109.720 174.525 ;
        RECT 109.890 174.325 110.220 174.525 ;
        RECT 107.585 174.135 107.815 174.185 ;
        RECT 107.585 173.505 107.925 174.135 ;
        RECT 108.095 173.335 108.345 174.135 ;
        RECT 108.535 173.985 109.760 174.155 ;
        RECT 108.535 173.505 108.865 173.985 ;
        RECT 109.035 173.335 109.260 173.795 ;
        RECT 109.430 173.505 109.760 173.985 ;
        RECT 110.390 174.115 110.560 174.745 ;
        RECT 110.745 174.325 111.095 174.575 ;
        RECT 111.265 174.255 111.785 174.795 ;
        RECT 110.390 173.505 110.890 174.115 ;
        RECT 111.955 174.085 112.475 174.625 ;
        RECT 114.240 174.200 114.590 175.450 ;
        RECT 118.205 174.745 118.435 175.885 ;
        RECT 118.605 174.735 118.935 175.715 ;
        RECT 119.105 174.745 119.315 175.885 ;
        RECT 119.545 174.795 120.755 175.885 ;
        RECT 120.930 175.450 126.275 175.885 ;
        RECT 111.265 173.335 112.475 174.085 ;
        RECT 116.070 173.880 116.410 174.710 ;
        RECT 118.185 174.325 118.515 174.575 ;
        RECT 112.650 173.335 117.995 173.880 ;
        RECT 118.205 173.335 118.435 174.155 ;
        RECT 118.685 174.135 118.935 174.735 ;
        RECT 119.545 174.255 120.065 174.795 ;
        RECT 118.605 173.505 118.935 174.135 ;
        RECT 119.105 173.335 119.315 174.155 ;
        RECT 120.235 174.085 120.755 174.625 ;
        RECT 122.520 174.200 122.870 175.450 ;
        RECT 126.445 174.795 127.655 175.885 ;
        RECT 119.545 173.335 120.755 174.085 ;
        RECT 124.350 173.880 124.690 174.710 ;
        RECT 126.445 174.255 126.965 174.795 ;
        RECT 127.135 174.085 127.655 174.625 ;
        RECT 120.930 173.335 126.275 173.880 ;
        RECT 126.445 173.335 127.655 174.085 ;
        RECT 14.580 173.165 127.740 173.335 ;
        RECT 14.665 172.415 15.875 173.165 ;
        RECT 14.665 171.875 15.185 172.415 ;
        RECT 16.965 172.395 20.475 173.165 ;
        RECT 20.650 172.620 25.995 173.165 ;
        RECT 26.170 172.620 31.515 173.165 ;
        RECT 31.690 172.620 37.035 173.165 ;
        RECT 15.355 171.705 15.875 172.245 ;
        RECT 14.665 170.615 15.875 171.705 ;
        RECT 16.965 171.705 18.655 172.225 ;
        RECT 18.825 171.875 20.475 172.395 ;
        RECT 16.965 170.615 20.475 171.705 ;
        RECT 22.240 171.050 22.590 172.300 ;
        RECT 24.070 171.790 24.410 172.620 ;
        RECT 27.760 171.050 28.110 172.300 ;
        RECT 29.590 171.790 29.930 172.620 ;
        RECT 33.280 171.050 33.630 172.300 ;
        RECT 35.110 171.790 35.450 172.620 ;
        RECT 37.205 172.440 37.495 173.165 ;
        RECT 37.665 172.365 38.005 172.995 ;
        RECT 38.175 172.365 38.425 173.165 ;
        RECT 38.615 172.515 38.945 172.995 ;
        RECT 39.115 172.705 39.340 173.165 ;
        RECT 39.510 172.515 39.840 172.995 ;
        RECT 20.650 170.615 25.995 171.050 ;
        RECT 26.170 170.615 31.515 171.050 ;
        RECT 31.690 170.615 37.035 171.050 ;
        RECT 37.205 170.615 37.495 171.780 ;
        RECT 37.665 171.755 37.840 172.365 ;
        RECT 38.615 172.345 39.840 172.515 ;
        RECT 40.470 172.385 40.970 172.995 ;
        RECT 41.805 172.490 42.065 172.995 ;
        RECT 42.245 172.785 42.575 173.165 ;
        RECT 42.755 172.615 42.925 172.995 ;
        RECT 38.010 172.005 38.705 172.175 ;
        RECT 38.535 171.755 38.705 172.005 ;
        RECT 38.880 171.975 39.300 172.175 ;
        RECT 39.470 171.975 39.800 172.175 ;
        RECT 39.970 171.975 40.300 172.175 ;
        RECT 40.470 171.755 40.640 172.385 ;
        RECT 40.825 171.925 41.175 172.175 ;
        RECT 37.665 170.785 38.005 171.755 ;
        RECT 38.175 170.615 38.345 171.755 ;
        RECT 38.535 171.585 40.970 171.755 ;
        RECT 38.615 170.615 38.865 171.415 ;
        RECT 39.510 170.785 39.840 171.585 ;
        RECT 40.140 170.615 40.470 171.415 ;
        RECT 40.640 170.785 40.970 171.585 ;
        RECT 41.805 171.690 41.975 172.490 ;
        RECT 42.260 172.445 42.925 172.615 ;
        RECT 42.260 172.190 42.430 172.445 ;
        RECT 44.105 172.365 44.445 172.995 ;
        RECT 44.615 172.365 44.865 173.165 ;
        RECT 45.055 172.515 45.385 172.995 ;
        RECT 45.555 172.705 45.780 173.165 ;
        RECT 45.950 172.515 46.280 172.995 ;
        RECT 42.145 171.860 42.430 172.190 ;
        RECT 42.665 171.895 42.995 172.265 ;
        RECT 42.260 171.715 42.430 171.860 ;
        RECT 44.105 171.755 44.280 172.365 ;
        RECT 45.055 172.345 46.280 172.515 ;
        RECT 46.910 172.385 47.410 172.995 ;
        RECT 44.450 172.005 45.145 172.175 ;
        RECT 44.975 171.755 45.145 172.005 ;
        RECT 45.320 171.975 45.740 172.175 ;
        RECT 45.910 171.975 46.240 172.175 ;
        RECT 46.410 171.975 46.740 172.175 ;
        RECT 46.910 171.755 47.080 172.385 ;
        RECT 47.785 172.365 48.125 172.995 ;
        RECT 48.295 172.365 48.545 173.165 ;
        RECT 48.735 172.515 49.065 172.995 ;
        RECT 49.235 172.705 49.460 173.165 ;
        RECT 49.630 172.515 49.960 172.995 ;
        RECT 47.265 171.925 47.615 172.175 ;
        RECT 47.785 171.755 47.960 172.365 ;
        RECT 48.735 172.345 49.960 172.515 ;
        RECT 50.590 172.385 51.090 172.995 ;
        RECT 48.130 172.005 48.825 172.175 ;
        RECT 48.655 171.755 48.825 172.005 ;
        RECT 49.000 171.975 49.420 172.175 ;
        RECT 49.590 171.975 49.920 172.175 ;
        RECT 50.090 171.975 50.420 172.175 ;
        RECT 50.590 171.755 50.760 172.385 ;
        RECT 51.465 172.365 51.805 172.995 ;
        RECT 51.975 172.365 52.225 173.165 ;
        RECT 52.415 172.515 52.745 172.995 ;
        RECT 52.915 172.705 53.140 173.165 ;
        RECT 53.310 172.515 53.640 172.995 ;
        RECT 50.945 171.925 51.295 172.175 ;
        RECT 51.465 171.755 51.640 172.365 ;
        RECT 52.415 172.345 53.640 172.515 ;
        RECT 54.270 172.385 54.770 172.995 ;
        RECT 55.145 172.415 56.355 173.165 ;
        RECT 51.810 172.005 52.505 172.175 ;
        RECT 52.335 171.755 52.505 172.005 ;
        RECT 52.680 171.975 53.100 172.175 ;
        RECT 53.270 171.975 53.600 172.175 ;
        RECT 53.770 171.975 54.100 172.175 ;
        RECT 54.270 171.755 54.440 172.385 ;
        RECT 54.625 171.925 54.975 172.175 ;
        RECT 41.805 170.785 42.075 171.690 ;
        RECT 42.260 171.545 42.925 171.715 ;
        RECT 42.245 170.615 42.575 171.375 ;
        RECT 42.755 170.785 42.925 171.545 ;
        RECT 44.105 170.785 44.445 171.755 ;
        RECT 44.615 170.615 44.785 171.755 ;
        RECT 44.975 171.585 47.410 171.755 ;
        RECT 45.055 170.615 45.305 171.415 ;
        RECT 45.950 170.785 46.280 171.585 ;
        RECT 46.580 170.615 46.910 171.415 ;
        RECT 47.080 170.785 47.410 171.585 ;
        RECT 47.785 170.785 48.125 171.755 ;
        RECT 48.295 170.615 48.465 171.755 ;
        RECT 48.655 171.585 51.090 171.755 ;
        RECT 48.735 170.615 48.985 171.415 ;
        RECT 49.630 170.785 49.960 171.585 ;
        RECT 50.260 170.615 50.590 171.415 ;
        RECT 50.760 170.785 51.090 171.585 ;
        RECT 51.465 170.785 51.805 171.755 ;
        RECT 51.975 170.615 52.145 171.755 ;
        RECT 52.335 171.585 54.770 171.755 ;
        RECT 52.415 170.615 52.665 171.415 ;
        RECT 53.310 170.785 53.640 171.585 ;
        RECT 53.940 170.615 54.270 171.415 ;
        RECT 54.440 170.785 54.770 171.585 ;
        RECT 55.145 171.705 55.665 172.245 ;
        RECT 55.835 171.875 56.355 172.415 ;
        RECT 56.525 172.395 60.035 173.165 ;
        RECT 56.525 171.705 58.215 172.225 ;
        RECT 58.385 171.875 60.035 172.395 ;
        RECT 60.265 172.345 60.475 173.165 ;
        RECT 60.645 172.365 60.975 172.995 ;
        RECT 60.645 171.765 60.895 172.365 ;
        RECT 61.145 172.345 61.375 173.165 ;
        RECT 61.675 172.615 61.845 172.995 ;
        RECT 62.025 172.785 62.355 173.165 ;
        RECT 61.675 172.445 62.340 172.615 ;
        RECT 62.535 172.490 62.795 172.995 ;
        RECT 61.065 171.925 61.395 172.175 ;
        RECT 61.605 171.895 61.935 172.265 ;
        RECT 62.170 172.190 62.340 172.445 ;
        RECT 62.170 171.860 62.455 172.190 ;
        RECT 55.145 170.615 56.355 171.705 ;
        RECT 56.525 170.615 60.035 171.705 ;
        RECT 60.265 170.615 60.475 171.755 ;
        RECT 60.645 170.785 60.975 171.765 ;
        RECT 61.145 170.615 61.375 171.755 ;
        RECT 62.170 171.715 62.340 171.860 ;
        RECT 61.675 171.545 62.340 171.715 ;
        RECT 62.625 171.690 62.795 172.490 ;
        RECT 62.965 172.440 63.255 173.165 ;
        RECT 63.885 172.395 65.555 173.165 ;
        RECT 65.730 172.620 71.075 173.165 ;
        RECT 71.250 172.620 76.595 173.165 ;
        RECT 76.770 172.620 82.115 173.165 ;
        RECT 61.675 170.785 61.845 171.545 ;
        RECT 62.025 170.615 62.355 171.375 ;
        RECT 62.525 170.785 62.795 171.690 ;
        RECT 62.965 170.615 63.255 171.780 ;
        RECT 63.885 171.705 64.635 172.225 ;
        RECT 64.805 171.875 65.555 172.395 ;
        RECT 63.885 170.615 65.555 171.705 ;
        RECT 67.320 171.050 67.670 172.300 ;
        RECT 69.150 171.790 69.490 172.620 ;
        RECT 72.840 171.050 73.190 172.300 ;
        RECT 74.670 171.790 75.010 172.620 ;
        RECT 78.360 171.050 78.710 172.300 ;
        RECT 80.190 171.790 80.530 172.620 ;
        RECT 82.375 172.515 82.545 172.995 ;
        RECT 82.725 172.685 82.965 173.165 ;
        RECT 83.215 172.515 83.385 172.995 ;
        RECT 83.555 172.685 83.885 173.165 ;
        RECT 84.055 172.515 84.225 172.995 ;
        RECT 82.375 172.345 83.010 172.515 ;
        RECT 83.215 172.345 84.225 172.515 ;
        RECT 84.395 172.365 84.725 173.165 ;
        RECT 85.160 172.535 85.445 172.995 ;
        RECT 85.615 172.705 85.885 173.165 ;
        RECT 85.160 172.365 86.115 172.535 ;
        RECT 82.840 172.175 83.010 172.345 ;
        RECT 83.725 172.315 84.225 172.345 ;
        RECT 82.290 171.935 82.670 172.175 ;
        RECT 82.840 172.005 83.340 172.175 ;
        RECT 82.840 171.765 83.010 172.005 ;
        RECT 83.730 171.805 84.225 172.315 ;
        RECT 82.295 171.595 83.010 171.765 ;
        RECT 83.215 171.635 84.225 171.805 ;
        RECT 65.730 170.615 71.075 171.050 ;
        RECT 71.250 170.615 76.595 171.050 ;
        RECT 76.770 170.615 82.115 171.050 ;
        RECT 82.295 170.785 82.625 171.595 ;
        RECT 82.795 170.615 83.035 171.415 ;
        RECT 83.215 170.785 83.385 171.635 ;
        RECT 83.555 170.615 83.885 171.415 ;
        RECT 84.055 170.785 84.225 171.635 ;
        RECT 84.395 170.615 84.725 171.765 ;
        RECT 85.045 171.635 85.735 172.195 ;
        RECT 85.905 171.465 86.115 172.365 ;
        RECT 85.160 171.245 86.115 171.465 ;
        RECT 86.285 172.195 86.685 172.995 ;
        RECT 86.875 172.535 87.155 172.995 ;
        RECT 87.675 172.705 88.000 173.165 ;
        RECT 86.875 172.365 88.000 172.535 ;
        RECT 88.170 172.425 88.555 172.995 ;
        RECT 88.725 172.440 89.015 173.165 ;
        RECT 87.550 172.255 88.000 172.365 ;
        RECT 86.285 171.635 87.380 172.195 ;
        RECT 87.550 171.925 88.105 172.255 ;
        RECT 85.160 170.785 85.445 171.245 ;
        RECT 85.615 170.615 85.885 171.075 ;
        RECT 86.285 170.785 86.685 171.635 ;
        RECT 87.550 171.465 88.000 171.925 ;
        RECT 88.275 171.755 88.555 172.425 ;
        RECT 89.685 172.345 89.915 173.165 ;
        RECT 90.085 172.365 90.415 172.995 ;
        RECT 89.665 171.925 89.995 172.175 ;
        RECT 86.875 171.245 88.000 171.465 ;
        RECT 86.875 170.785 87.155 171.245 ;
        RECT 87.675 170.615 88.000 171.075 ;
        RECT 88.170 170.785 88.555 171.755 ;
        RECT 88.725 170.615 89.015 171.780 ;
        RECT 90.165 171.765 90.415 172.365 ;
        RECT 90.585 172.345 90.795 173.165 ;
        RECT 91.030 172.455 91.285 172.985 ;
        RECT 91.455 172.705 91.760 173.165 ;
        RECT 92.005 172.785 93.075 172.955 ;
        RECT 89.685 170.615 89.915 171.755 ;
        RECT 90.085 170.785 90.415 171.765 ;
        RECT 91.030 171.805 91.240 172.455 ;
        RECT 92.005 172.430 92.325 172.785 ;
        RECT 92.000 172.255 92.325 172.430 ;
        RECT 91.410 171.955 92.325 172.255 ;
        RECT 92.495 172.215 92.735 172.615 ;
        RECT 92.905 172.555 93.075 172.785 ;
        RECT 93.245 172.725 93.435 173.165 ;
        RECT 93.605 172.715 94.555 172.995 ;
        RECT 94.775 172.805 95.125 172.975 ;
        RECT 92.905 172.385 93.435 172.555 ;
        RECT 91.410 171.925 92.150 171.955 ;
        RECT 90.585 170.615 90.795 171.755 ;
        RECT 91.030 170.925 91.285 171.805 ;
        RECT 91.455 170.615 91.760 171.755 ;
        RECT 91.980 171.335 92.150 171.925 ;
        RECT 92.495 171.845 93.035 172.215 ;
        RECT 93.215 172.105 93.435 172.385 ;
        RECT 93.605 171.935 93.775 172.715 ;
        RECT 93.370 171.765 93.775 171.935 ;
        RECT 93.945 171.925 94.295 172.545 ;
        RECT 93.370 171.675 93.540 171.765 ;
        RECT 94.465 171.755 94.675 172.545 ;
        RECT 92.320 171.505 93.540 171.675 ;
        RECT 94.000 171.595 94.675 171.755 ;
        RECT 91.980 171.165 92.780 171.335 ;
        RECT 92.100 170.615 92.430 170.995 ;
        RECT 92.610 170.875 92.780 171.165 ;
        RECT 93.370 171.125 93.540 171.505 ;
        RECT 93.710 171.585 94.675 171.595 ;
        RECT 94.865 172.415 95.125 172.805 ;
        RECT 95.335 172.705 95.665 173.165 ;
        RECT 96.540 172.775 97.395 172.945 ;
        RECT 97.600 172.775 98.095 172.945 ;
        RECT 98.265 172.805 98.595 173.165 ;
        RECT 94.865 171.725 95.035 172.415 ;
        RECT 95.205 172.065 95.375 172.245 ;
        RECT 95.545 172.235 96.335 172.485 ;
        RECT 96.540 172.065 96.710 172.775 ;
        RECT 96.880 172.265 97.235 172.485 ;
        RECT 95.205 171.895 96.895 172.065 ;
        RECT 93.710 171.295 94.170 171.585 ;
        RECT 94.865 171.555 96.365 171.725 ;
        RECT 94.865 171.415 95.035 171.555 ;
        RECT 94.475 171.245 95.035 171.415 ;
        RECT 92.950 170.615 93.200 171.075 ;
        RECT 93.370 170.785 94.240 171.125 ;
        RECT 94.475 170.785 94.645 171.245 ;
        RECT 95.480 171.215 96.555 171.385 ;
        RECT 94.815 170.615 95.185 171.075 ;
        RECT 95.480 170.875 95.650 171.215 ;
        RECT 95.820 170.615 96.150 171.045 ;
        RECT 96.385 170.875 96.555 171.215 ;
        RECT 96.725 171.115 96.895 171.895 ;
        RECT 97.065 171.675 97.235 172.265 ;
        RECT 97.405 171.865 97.755 172.485 ;
        RECT 97.065 171.285 97.530 171.675 ;
        RECT 97.925 171.415 98.095 172.775 ;
        RECT 98.265 171.585 98.725 172.635 ;
        RECT 97.700 171.245 98.095 171.415 ;
        RECT 97.700 171.115 97.870 171.245 ;
        RECT 96.725 170.785 97.405 171.115 ;
        RECT 97.620 170.785 97.870 171.115 ;
        RECT 98.040 170.615 98.290 171.075 ;
        RECT 98.460 170.800 98.785 171.585 ;
        RECT 98.955 170.785 99.125 172.905 ;
        RECT 99.295 172.785 99.625 173.165 ;
        RECT 99.795 172.615 100.050 172.905 ;
        RECT 101.150 172.620 106.495 173.165 ;
        RECT 99.300 172.445 100.050 172.615 ;
        RECT 99.300 171.455 99.530 172.445 ;
        RECT 99.700 171.625 100.050 172.275 ;
        RECT 99.300 171.285 100.050 171.455 ;
        RECT 99.295 170.615 99.625 171.115 ;
        RECT 99.795 170.785 100.050 171.285 ;
        RECT 102.740 171.050 103.090 172.300 ;
        RECT 104.570 171.790 104.910 172.620 ;
        RECT 106.725 172.345 106.935 173.165 ;
        RECT 107.105 172.365 107.435 172.995 ;
        RECT 107.105 171.765 107.355 172.365 ;
        RECT 107.605 172.345 107.835 173.165 ;
        RECT 108.250 172.385 108.750 172.995 ;
        RECT 107.525 171.925 107.855 172.175 ;
        RECT 108.045 171.925 108.395 172.175 ;
        RECT 101.150 170.615 106.495 171.050 ;
        RECT 106.725 170.615 106.935 171.755 ;
        RECT 107.105 170.785 107.435 171.765 ;
        RECT 108.580 171.755 108.750 172.385 ;
        RECT 109.380 172.515 109.710 172.995 ;
        RECT 109.880 172.705 110.105 173.165 ;
        RECT 110.275 172.515 110.605 172.995 ;
        RECT 109.380 172.345 110.605 172.515 ;
        RECT 110.795 172.365 111.045 173.165 ;
        RECT 111.215 172.365 111.555 172.995 ;
        RECT 111.725 172.415 112.935 173.165 ;
        RECT 108.920 171.975 109.250 172.175 ;
        RECT 109.420 171.975 109.750 172.175 ;
        RECT 109.920 171.975 110.340 172.175 ;
        RECT 110.515 172.005 111.210 172.175 ;
        RECT 110.515 171.755 110.685 172.005 ;
        RECT 111.380 171.755 111.555 172.365 ;
        RECT 107.605 170.615 107.835 171.755 ;
        RECT 108.250 171.585 110.685 171.755 ;
        RECT 108.250 170.785 108.580 171.585 ;
        RECT 108.750 170.615 109.080 171.415 ;
        RECT 109.380 170.785 109.710 171.585 ;
        RECT 110.355 170.615 110.605 171.415 ;
        RECT 110.875 170.615 111.045 171.755 ;
        RECT 111.215 170.785 111.555 171.755 ;
        RECT 111.725 171.705 112.245 172.245 ;
        RECT 112.415 171.875 112.935 172.415 ;
        RECT 113.145 172.345 113.375 173.165 ;
        RECT 113.545 172.365 113.875 172.995 ;
        RECT 113.125 171.925 113.455 172.175 ;
        RECT 113.625 171.765 113.875 172.365 ;
        RECT 114.045 172.345 114.255 173.165 ;
        RECT 114.485 172.440 114.775 173.165 ;
        RECT 115.870 172.455 116.125 172.985 ;
        RECT 116.295 172.705 116.600 173.165 ;
        RECT 116.845 172.785 117.915 172.955 ;
        RECT 115.870 171.805 116.080 172.455 ;
        RECT 116.845 172.430 117.165 172.785 ;
        RECT 116.840 172.255 117.165 172.430 ;
        RECT 116.250 171.955 117.165 172.255 ;
        RECT 117.335 172.215 117.575 172.615 ;
        RECT 117.745 172.555 117.915 172.785 ;
        RECT 118.085 172.725 118.275 173.165 ;
        RECT 118.445 172.715 119.395 172.995 ;
        RECT 119.615 172.805 119.965 172.975 ;
        RECT 117.745 172.385 118.275 172.555 ;
        RECT 116.250 171.925 116.990 171.955 ;
        RECT 111.725 170.615 112.935 171.705 ;
        RECT 113.145 170.615 113.375 171.755 ;
        RECT 113.545 170.785 113.875 171.765 ;
        RECT 114.045 170.615 114.255 171.755 ;
        RECT 114.485 170.615 114.775 171.780 ;
        RECT 115.870 170.925 116.125 171.805 ;
        RECT 116.295 170.615 116.600 171.755 ;
        RECT 116.820 171.335 116.990 171.925 ;
        RECT 117.335 171.845 117.875 172.215 ;
        RECT 118.055 172.105 118.275 172.385 ;
        RECT 118.445 171.935 118.615 172.715 ;
        RECT 118.210 171.765 118.615 171.935 ;
        RECT 118.785 171.925 119.135 172.545 ;
        RECT 118.210 171.675 118.380 171.765 ;
        RECT 119.305 171.755 119.515 172.545 ;
        RECT 117.160 171.505 118.380 171.675 ;
        RECT 118.840 171.595 119.515 171.755 ;
        RECT 116.820 171.165 117.620 171.335 ;
        RECT 116.940 170.615 117.270 170.995 ;
        RECT 117.450 170.875 117.620 171.165 ;
        RECT 118.210 171.125 118.380 171.505 ;
        RECT 118.550 171.585 119.515 171.595 ;
        RECT 119.705 172.415 119.965 172.805 ;
        RECT 120.175 172.705 120.505 173.165 ;
        RECT 121.380 172.775 122.235 172.945 ;
        RECT 122.440 172.775 122.935 172.945 ;
        RECT 123.105 172.805 123.435 173.165 ;
        RECT 119.705 171.725 119.875 172.415 ;
        RECT 120.045 172.065 120.215 172.245 ;
        RECT 120.385 172.235 121.175 172.485 ;
        RECT 121.380 172.065 121.550 172.775 ;
        RECT 121.720 172.265 122.075 172.485 ;
        RECT 120.045 171.895 121.735 172.065 ;
        RECT 118.550 171.295 119.010 171.585 ;
        RECT 119.705 171.555 121.205 171.725 ;
        RECT 119.705 171.415 119.875 171.555 ;
        RECT 119.315 171.245 119.875 171.415 ;
        RECT 117.790 170.615 118.040 171.075 ;
        RECT 118.210 170.785 119.080 171.125 ;
        RECT 119.315 170.785 119.485 171.245 ;
        RECT 120.320 171.215 121.395 171.385 ;
        RECT 119.655 170.615 120.025 171.075 ;
        RECT 120.320 170.875 120.490 171.215 ;
        RECT 120.660 170.615 120.990 171.045 ;
        RECT 121.225 170.875 121.395 171.215 ;
        RECT 121.565 171.115 121.735 171.895 ;
        RECT 121.905 171.675 122.075 172.265 ;
        RECT 122.245 171.865 122.595 172.485 ;
        RECT 121.905 171.285 122.370 171.675 ;
        RECT 122.765 171.415 122.935 172.775 ;
        RECT 123.105 171.585 123.565 172.635 ;
        RECT 122.540 171.245 122.935 171.415 ;
        RECT 122.540 171.115 122.710 171.245 ;
        RECT 121.565 170.785 122.245 171.115 ;
        RECT 122.460 170.785 122.710 171.115 ;
        RECT 122.880 170.615 123.130 171.075 ;
        RECT 123.300 170.800 123.625 171.585 ;
        RECT 123.795 170.785 123.965 172.905 ;
        RECT 124.135 172.785 124.465 173.165 ;
        RECT 124.635 172.615 124.890 172.905 ;
        RECT 124.140 172.445 124.890 172.615 ;
        RECT 124.140 171.455 124.370 172.445 ;
        RECT 125.065 172.415 126.275 173.165 ;
        RECT 126.445 172.415 127.655 173.165 ;
        RECT 124.540 171.625 124.890 172.275 ;
        RECT 125.065 171.705 125.585 172.245 ;
        RECT 125.755 171.875 126.275 172.415 ;
        RECT 126.445 171.705 126.965 172.245 ;
        RECT 127.135 171.875 127.655 172.415 ;
        RECT 124.140 171.285 124.890 171.455 ;
        RECT 124.135 170.615 124.465 171.115 ;
        RECT 124.635 170.785 124.890 171.285 ;
        RECT 125.065 170.615 126.275 171.705 ;
        RECT 126.445 170.615 127.655 171.705 ;
        RECT 14.580 170.445 127.740 170.615 ;
        RECT 14.665 169.355 15.875 170.445 ;
        RECT 14.665 168.645 15.185 169.185 ;
        RECT 15.355 168.815 15.875 169.355 ;
        RECT 16.045 169.355 18.635 170.445 ;
        RECT 18.810 170.010 24.155 170.445 ;
        RECT 16.045 168.835 17.255 169.355 ;
        RECT 17.425 168.665 18.635 169.185 ;
        RECT 20.400 168.760 20.750 170.010 ;
        RECT 24.325 169.280 24.615 170.445 ;
        RECT 25.245 169.355 26.915 170.445 ;
        RECT 14.665 167.895 15.875 168.645 ;
        RECT 16.045 167.895 18.635 168.665 ;
        RECT 22.230 168.440 22.570 169.270 ;
        RECT 25.245 168.835 25.995 169.355 ;
        RECT 27.125 169.305 27.355 170.445 ;
        RECT 27.525 169.295 27.855 170.275 ;
        RECT 28.025 169.305 28.235 170.445 ;
        RECT 28.925 169.355 32.435 170.445 ;
        RECT 26.165 168.665 26.915 169.185 ;
        RECT 27.105 168.885 27.435 169.135 ;
        RECT 18.810 167.895 24.155 168.440 ;
        RECT 24.325 167.895 24.615 168.620 ;
        RECT 25.245 167.895 26.915 168.665 ;
        RECT 27.125 167.895 27.355 168.715 ;
        RECT 27.605 168.695 27.855 169.295 ;
        RECT 28.925 168.835 30.615 169.355 ;
        RECT 32.665 169.305 32.875 170.445 ;
        RECT 33.045 169.295 33.375 170.275 ;
        RECT 33.545 169.305 33.775 170.445 ;
        RECT 33.985 169.355 35.195 170.445 ;
        RECT 35.455 169.700 35.725 170.445 ;
        RECT 36.355 170.440 42.630 170.445 ;
        RECT 35.895 169.530 36.185 170.270 ;
        RECT 36.355 169.715 36.610 170.440 ;
        RECT 36.795 169.545 37.055 170.270 ;
        RECT 37.225 169.715 37.470 170.440 ;
        RECT 37.655 169.545 37.915 170.270 ;
        RECT 38.085 169.715 38.330 170.440 ;
        RECT 38.515 169.545 38.775 170.270 ;
        RECT 38.945 169.715 39.190 170.440 ;
        RECT 39.360 169.545 39.620 170.270 ;
        RECT 39.790 169.715 40.050 170.440 ;
        RECT 40.220 169.545 40.480 170.270 ;
        RECT 40.650 169.715 40.910 170.440 ;
        RECT 41.080 169.545 41.340 170.270 ;
        RECT 41.510 169.715 41.770 170.440 ;
        RECT 41.940 169.545 42.200 170.270 ;
        RECT 42.370 169.645 42.630 170.440 ;
        RECT 36.795 169.530 42.200 169.545 ;
        RECT 27.525 168.065 27.855 168.695 ;
        RECT 28.025 167.895 28.235 168.715 ;
        RECT 30.785 168.665 32.435 169.185 ;
        RECT 28.925 167.895 32.435 168.665 ;
        RECT 32.665 167.895 32.875 168.715 ;
        RECT 33.045 168.695 33.295 169.295 ;
        RECT 33.465 168.885 33.795 169.135 ;
        RECT 33.985 168.815 34.505 169.355 ;
        RECT 35.455 169.305 42.200 169.530 ;
        RECT 33.045 168.065 33.375 168.695 ;
        RECT 33.545 167.895 33.775 168.715 ;
        RECT 34.675 168.645 35.195 169.185 ;
        RECT 33.985 167.895 35.195 168.645 ;
        RECT 35.455 168.715 36.620 169.305 ;
        RECT 42.800 169.135 43.050 170.270 ;
        RECT 43.230 169.635 43.490 170.445 ;
        RECT 43.665 169.135 43.910 170.275 ;
        RECT 44.090 169.635 44.385 170.445 ;
        RECT 44.570 170.010 49.915 170.445 ;
        RECT 36.790 168.885 43.910 169.135 ;
        RECT 35.455 168.545 42.200 168.715 ;
        RECT 35.455 167.895 35.755 168.375 ;
        RECT 35.925 168.090 36.185 168.545 ;
        RECT 36.355 167.895 36.615 168.375 ;
        RECT 36.795 168.090 37.055 168.545 ;
        RECT 37.225 167.895 37.475 168.375 ;
        RECT 37.655 168.090 37.915 168.545 ;
        RECT 38.085 167.895 38.335 168.375 ;
        RECT 38.515 168.090 38.775 168.545 ;
        RECT 38.945 167.895 39.190 168.375 ;
        RECT 39.360 168.090 39.635 168.545 ;
        RECT 39.805 167.895 40.050 168.375 ;
        RECT 40.220 168.090 40.480 168.545 ;
        RECT 40.650 167.895 40.910 168.375 ;
        RECT 41.080 168.090 41.340 168.545 ;
        RECT 41.510 167.895 41.770 168.375 ;
        RECT 41.940 168.090 42.200 168.545 ;
        RECT 42.370 167.895 42.630 168.455 ;
        RECT 42.800 168.075 43.050 168.885 ;
        RECT 43.230 167.895 43.490 168.420 ;
        RECT 43.660 168.075 43.910 168.885 ;
        RECT 44.080 168.575 44.395 169.135 ;
        RECT 46.160 168.760 46.510 170.010 ;
        RECT 50.085 169.280 50.375 170.445 ;
        RECT 50.545 169.355 51.755 170.445 ;
        RECT 51.930 170.010 57.275 170.445 ;
        RECT 57.450 170.010 62.795 170.445 ;
        RECT 62.970 170.010 68.315 170.445 ;
        RECT 47.990 168.440 48.330 169.270 ;
        RECT 50.545 168.815 51.065 169.355 ;
        RECT 51.235 168.645 51.755 169.185 ;
        RECT 53.520 168.760 53.870 170.010 ;
        RECT 44.090 167.895 44.395 168.405 ;
        RECT 44.570 167.895 49.915 168.440 ;
        RECT 50.085 167.895 50.375 168.620 ;
        RECT 50.545 167.895 51.755 168.645 ;
        RECT 55.350 168.440 55.690 169.270 ;
        RECT 59.040 168.760 59.390 170.010 ;
        RECT 60.870 168.440 61.210 169.270 ;
        RECT 64.560 168.760 64.910 170.010 ;
        RECT 68.490 169.295 68.750 170.445 ;
        RECT 68.925 169.370 69.180 170.275 ;
        RECT 69.350 169.685 69.680 170.445 ;
        RECT 69.895 169.515 70.065 170.275 ;
        RECT 66.390 168.440 66.730 169.270 ;
        RECT 51.930 167.895 57.275 168.440 ;
        RECT 57.450 167.895 62.795 168.440 ;
        RECT 62.970 167.895 68.315 168.440 ;
        RECT 68.490 167.895 68.750 168.735 ;
        RECT 68.925 168.640 69.095 169.370 ;
        RECT 69.350 169.345 70.065 169.515 ;
        RECT 69.350 169.135 69.520 169.345 ;
        RECT 70.330 169.295 70.590 170.445 ;
        RECT 70.765 169.370 71.020 170.275 ;
        RECT 71.190 169.685 71.520 170.445 ;
        RECT 71.735 169.515 71.905 170.275 ;
        RECT 69.265 168.805 69.520 169.135 ;
        RECT 68.925 168.065 69.180 168.640 ;
        RECT 69.350 168.615 69.520 168.805 ;
        RECT 69.800 168.795 70.155 169.165 ;
        RECT 69.350 168.445 70.065 168.615 ;
        RECT 69.350 167.895 69.680 168.275 ;
        RECT 69.895 168.065 70.065 168.445 ;
        RECT 70.330 167.895 70.590 168.735 ;
        RECT 70.765 168.640 70.935 169.370 ;
        RECT 71.190 169.345 71.905 169.515 ;
        RECT 72.165 169.355 75.675 170.445 ;
        RECT 71.190 169.135 71.360 169.345 ;
        RECT 71.105 168.805 71.360 169.135 ;
        RECT 70.765 168.065 71.020 168.640 ;
        RECT 71.190 168.615 71.360 168.805 ;
        RECT 71.640 168.795 71.995 169.165 ;
        RECT 72.165 168.835 73.855 169.355 ;
        RECT 75.845 169.280 76.135 170.445 ;
        RECT 76.305 169.685 76.820 170.095 ;
        RECT 77.055 169.685 77.225 170.445 ;
        RECT 77.395 170.105 79.425 170.275 ;
        RECT 74.025 168.665 75.675 169.185 ;
        RECT 76.305 168.875 76.645 169.685 ;
        RECT 77.395 169.440 77.565 170.105 ;
        RECT 77.960 169.765 79.085 169.935 ;
        RECT 76.815 169.250 77.565 169.440 ;
        RECT 77.735 169.425 78.745 169.595 ;
        RECT 76.305 168.705 77.535 168.875 ;
        RECT 71.190 168.445 71.905 168.615 ;
        RECT 71.190 167.895 71.520 168.275 ;
        RECT 71.735 168.065 71.905 168.445 ;
        RECT 72.165 167.895 75.675 168.665 ;
        RECT 75.845 167.895 76.135 168.620 ;
        RECT 76.580 168.100 76.825 168.705 ;
        RECT 77.045 167.895 77.555 168.430 ;
        RECT 77.735 168.065 77.925 169.425 ;
        RECT 78.095 168.405 78.370 169.225 ;
        RECT 78.575 168.625 78.745 169.425 ;
        RECT 78.915 168.635 79.085 169.765 ;
        RECT 79.255 169.135 79.425 170.105 ;
        RECT 79.595 169.305 79.765 170.445 ;
        RECT 79.935 169.305 80.270 170.275 ;
        RECT 79.255 168.805 79.450 169.135 ;
        RECT 79.675 168.805 79.930 169.135 ;
        RECT 79.675 168.635 79.845 168.805 ;
        RECT 80.100 168.635 80.270 169.305 ;
        RECT 80.820 169.465 81.075 170.135 ;
        RECT 81.255 169.645 81.540 170.445 ;
        RECT 81.720 169.725 82.050 170.235 ;
        RECT 80.820 168.745 81.000 169.465 ;
        RECT 81.720 169.135 81.970 169.725 ;
        RECT 82.320 169.575 82.490 170.185 ;
        RECT 82.660 169.755 82.990 170.445 ;
        RECT 83.220 169.895 83.460 170.185 ;
        RECT 83.660 170.065 84.080 170.445 ;
        RECT 84.260 169.975 84.890 170.225 ;
        RECT 85.360 170.065 85.690 170.445 ;
        RECT 84.260 169.895 84.430 169.975 ;
        RECT 85.860 169.895 86.030 170.185 ;
        RECT 86.210 170.065 86.590 170.445 ;
        RECT 86.830 170.060 87.660 170.230 ;
        RECT 83.220 169.725 84.430 169.895 ;
        RECT 81.170 168.805 81.970 169.135 ;
        RECT 78.915 168.465 79.845 168.635 ;
        RECT 78.915 168.430 79.090 168.465 ;
        RECT 78.095 168.235 78.375 168.405 ;
        RECT 78.095 168.065 78.370 168.235 ;
        RECT 78.560 168.065 79.090 168.430 ;
        RECT 79.515 167.895 79.845 168.295 ;
        RECT 80.015 168.065 80.270 168.635 ;
        RECT 80.735 168.605 81.000 168.745 ;
        RECT 80.735 168.575 81.075 168.605 ;
        RECT 80.820 168.075 81.075 168.575 ;
        RECT 81.255 167.895 81.540 168.355 ;
        RECT 81.720 168.155 81.970 168.805 ;
        RECT 82.170 169.555 82.490 169.575 ;
        RECT 82.170 169.385 84.090 169.555 ;
        RECT 82.170 168.490 82.360 169.385 ;
        RECT 84.260 169.215 84.430 169.725 ;
        RECT 84.600 169.465 85.120 169.775 ;
        RECT 82.530 169.045 84.430 169.215 ;
        RECT 82.530 168.985 82.860 169.045 ;
        RECT 83.010 168.815 83.340 168.875 ;
        RECT 82.680 168.545 83.340 168.815 ;
        RECT 82.170 168.160 82.490 168.490 ;
        RECT 82.670 167.895 83.330 168.375 ;
        RECT 83.530 168.285 83.700 169.045 ;
        RECT 84.600 168.875 84.780 169.285 ;
        RECT 83.870 168.705 84.200 168.825 ;
        RECT 84.950 168.705 85.120 169.465 ;
        RECT 83.870 168.535 85.120 168.705 ;
        RECT 85.290 169.645 86.660 169.895 ;
        RECT 85.290 168.875 85.480 169.645 ;
        RECT 86.410 169.385 86.660 169.645 ;
        RECT 85.650 169.215 85.900 169.375 ;
        RECT 86.830 169.215 87.000 170.060 ;
        RECT 87.895 169.775 88.065 170.275 ;
        RECT 88.235 169.945 88.565 170.445 ;
        RECT 87.170 169.385 87.670 169.765 ;
        RECT 87.895 169.605 88.590 169.775 ;
        RECT 85.650 169.045 87.000 169.215 ;
        RECT 86.580 169.005 87.000 169.045 ;
        RECT 85.290 168.535 85.710 168.875 ;
        RECT 86.000 168.545 86.410 168.875 ;
        RECT 83.530 168.115 84.380 168.285 ;
        RECT 84.940 167.895 85.260 168.355 ;
        RECT 85.460 168.105 85.710 168.535 ;
        RECT 86.000 167.895 86.410 168.335 ;
        RECT 86.580 168.275 86.750 169.005 ;
        RECT 86.920 168.455 87.270 168.825 ;
        RECT 87.450 168.515 87.670 169.385 ;
        RECT 87.840 168.815 88.250 169.435 ;
        RECT 88.420 168.635 88.590 169.605 ;
        RECT 87.895 168.445 88.590 168.635 ;
        RECT 86.580 168.075 87.595 168.275 ;
        RECT 87.895 168.115 88.065 168.445 ;
        RECT 88.235 167.895 88.565 168.275 ;
        RECT 88.780 168.155 89.005 170.275 ;
        RECT 89.175 169.945 89.505 170.445 ;
        RECT 89.675 169.775 89.845 170.275 ;
        RECT 89.180 169.605 89.845 169.775 ;
        RECT 89.180 168.615 89.410 169.605 ;
        RECT 89.580 168.785 89.930 169.435 ;
        RECT 90.105 169.355 91.315 170.445 ;
        RECT 91.485 169.685 92.000 170.095 ;
        RECT 92.235 169.685 92.405 170.445 ;
        RECT 92.575 170.105 94.605 170.275 ;
        RECT 90.105 168.815 90.625 169.355 ;
        RECT 90.795 168.645 91.315 169.185 ;
        RECT 91.485 168.875 91.825 169.685 ;
        RECT 92.575 169.440 92.745 170.105 ;
        RECT 93.140 169.765 94.265 169.935 ;
        RECT 91.995 169.250 92.745 169.440 ;
        RECT 92.915 169.425 93.925 169.595 ;
        RECT 91.485 168.705 92.715 168.875 ;
        RECT 89.180 168.445 89.845 168.615 ;
        RECT 89.175 167.895 89.505 168.275 ;
        RECT 89.675 168.155 89.845 168.445 ;
        RECT 90.105 167.895 91.315 168.645 ;
        RECT 91.760 168.100 92.005 168.705 ;
        RECT 92.225 167.895 92.735 168.430 ;
        RECT 92.915 168.065 93.105 169.425 ;
        RECT 93.275 169.085 93.550 169.225 ;
        RECT 93.275 168.915 93.555 169.085 ;
        RECT 93.275 168.065 93.550 168.915 ;
        RECT 93.755 168.625 93.925 169.425 ;
        RECT 94.095 168.635 94.265 169.765 ;
        RECT 94.435 169.135 94.605 170.105 ;
        RECT 94.775 169.305 94.945 170.445 ;
        RECT 95.115 169.305 95.450 170.275 ;
        RECT 96.175 169.515 96.345 170.275 ;
        RECT 96.525 169.685 96.855 170.445 ;
        RECT 96.175 169.345 96.840 169.515 ;
        RECT 97.025 169.370 97.295 170.275 ;
        RECT 94.435 168.805 94.630 169.135 ;
        RECT 94.855 168.805 95.110 169.135 ;
        RECT 94.855 168.635 95.025 168.805 ;
        RECT 95.280 168.635 95.450 169.305 ;
        RECT 96.670 169.200 96.840 169.345 ;
        RECT 96.105 168.795 96.435 169.165 ;
        RECT 96.670 168.870 96.955 169.200 ;
        RECT 94.095 168.465 95.025 168.635 ;
        RECT 94.095 168.430 94.270 168.465 ;
        RECT 93.740 168.065 94.270 168.430 ;
        RECT 94.695 167.895 95.025 168.295 ;
        RECT 95.195 168.065 95.450 168.635 ;
        RECT 96.670 168.615 96.840 168.870 ;
        RECT 96.175 168.445 96.840 168.615 ;
        RECT 97.125 168.570 97.295 169.370 ;
        RECT 97.925 169.355 101.435 170.445 ;
        RECT 97.925 168.835 99.615 169.355 ;
        RECT 101.605 169.280 101.895 170.445 ;
        RECT 102.990 169.255 103.245 170.135 ;
        RECT 103.415 169.305 103.720 170.445 ;
        RECT 104.060 170.065 104.390 170.445 ;
        RECT 104.570 169.895 104.740 170.185 ;
        RECT 104.910 169.985 105.160 170.445 ;
        RECT 103.940 169.725 104.740 169.895 ;
        RECT 105.330 169.935 106.200 170.275 ;
        RECT 99.785 168.665 101.435 169.185 ;
        RECT 96.175 168.065 96.345 168.445 ;
        RECT 96.525 167.895 96.855 168.275 ;
        RECT 97.035 168.065 97.295 168.570 ;
        RECT 97.925 167.895 101.435 168.665 ;
        RECT 101.605 167.895 101.895 168.620 ;
        RECT 102.990 168.605 103.200 169.255 ;
        RECT 103.940 169.135 104.110 169.725 ;
        RECT 105.330 169.555 105.500 169.935 ;
        RECT 106.435 169.815 106.605 170.275 ;
        RECT 106.775 169.985 107.145 170.445 ;
        RECT 107.440 169.845 107.610 170.185 ;
        RECT 107.780 170.015 108.110 170.445 ;
        RECT 108.345 169.845 108.515 170.185 ;
        RECT 104.280 169.385 105.500 169.555 ;
        RECT 105.670 169.475 106.130 169.765 ;
        RECT 106.435 169.645 106.995 169.815 ;
        RECT 107.440 169.675 108.515 169.845 ;
        RECT 108.685 169.945 109.365 170.275 ;
        RECT 109.580 169.945 109.830 170.275 ;
        RECT 110.000 169.985 110.250 170.445 ;
        RECT 106.825 169.505 106.995 169.645 ;
        RECT 105.670 169.465 106.635 169.475 ;
        RECT 105.330 169.295 105.500 169.385 ;
        RECT 105.960 169.305 106.635 169.465 ;
        RECT 103.370 169.105 104.110 169.135 ;
        RECT 103.370 168.805 104.285 169.105 ;
        RECT 103.960 168.630 104.285 168.805 ;
        RECT 102.990 168.075 103.245 168.605 ;
        RECT 103.415 167.895 103.720 168.355 ;
        RECT 103.965 168.275 104.285 168.630 ;
        RECT 104.455 168.845 104.995 169.215 ;
        RECT 105.330 169.125 105.735 169.295 ;
        RECT 104.455 168.445 104.695 168.845 ;
        RECT 105.175 168.675 105.395 168.955 ;
        RECT 104.865 168.505 105.395 168.675 ;
        RECT 104.865 168.275 105.035 168.505 ;
        RECT 105.565 168.345 105.735 169.125 ;
        RECT 105.905 168.515 106.255 169.135 ;
        RECT 106.425 168.515 106.635 169.305 ;
        RECT 106.825 169.335 108.325 169.505 ;
        RECT 106.825 168.645 106.995 169.335 ;
        RECT 108.685 169.165 108.855 169.945 ;
        RECT 109.660 169.815 109.830 169.945 ;
        RECT 107.165 168.995 108.855 169.165 ;
        RECT 109.025 169.385 109.490 169.775 ;
        RECT 109.660 169.645 110.055 169.815 ;
        RECT 107.165 168.815 107.335 168.995 ;
        RECT 103.965 168.105 105.035 168.275 ;
        RECT 105.205 167.895 105.395 168.335 ;
        RECT 105.565 168.065 106.515 168.345 ;
        RECT 106.825 168.255 107.085 168.645 ;
        RECT 107.505 168.575 108.295 168.825 ;
        RECT 106.735 168.085 107.085 168.255 ;
        RECT 107.295 167.895 107.625 168.355 ;
        RECT 108.500 168.285 108.670 168.995 ;
        RECT 109.025 168.795 109.195 169.385 ;
        RECT 108.840 168.575 109.195 168.795 ;
        RECT 109.365 168.575 109.715 169.195 ;
        RECT 109.885 168.285 110.055 169.645 ;
        RECT 110.420 169.475 110.745 170.260 ;
        RECT 110.225 168.425 110.685 169.475 ;
        RECT 108.500 168.115 109.355 168.285 ;
        RECT 109.560 168.115 110.055 168.285 ;
        RECT 110.225 167.895 110.555 168.255 ;
        RECT 110.915 168.155 111.085 170.275 ;
        RECT 111.255 169.945 111.585 170.445 ;
        RECT 111.755 169.775 112.010 170.275 ;
        RECT 111.260 169.605 112.010 169.775 ;
        RECT 111.260 168.615 111.490 169.605 ;
        RECT 111.660 168.785 112.010 169.435 ;
        RECT 112.650 169.305 112.985 170.275 ;
        RECT 113.155 169.305 113.325 170.445 ;
        RECT 113.495 170.105 115.525 170.275 ;
        RECT 112.650 168.635 112.820 169.305 ;
        RECT 113.495 169.135 113.665 170.105 ;
        RECT 112.990 168.805 113.245 169.135 ;
        RECT 113.470 168.805 113.665 169.135 ;
        RECT 113.835 169.765 114.960 169.935 ;
        RECT 113.075 168.635 113.245 168.805 ;
        RECT 113.835 168.635 114.005 169.765 ;
        RECT 111.260 168.445 112.010 168.615 ;
        RECT 111.255 167.895 111.585 168.275 ;
        RECT 111.755 168.155 112.010 168.445 ;
        RECT 112.650 168.065 112.905 168.635 ;
        RECT 113.075 168.465 114.005 168.635 ;
        RECT 114.175 169.425 115.185 169.595 ;
        RECT 114.175 168.625 114.345 169.425 ;
        RECT 114.550 169.085 114.825 169.225 ;
        RECT 114.545 168.915 114.825 169.085 ;
        RECT 113.830 168.430 114.005 168.465 ;
        RECT 113.075 167.895 113.405 168.295 ;
        RECT 113.830 168.065 114.360 168.430 ;
        RECT 114.550 168.065 114.825 168.915 ;
        RECT 114.995 168.065 115.185 169.425 ;
        RECT 115.355 169.440 115.525 170.105 ;
        RECT 115.695 169.685 115.865 170.445 ;
        RECT 116.100 169.685 116.615 170.095 ;
        RECT 115.355 169.250 116.105 169.440 ;
        RECT 116.275 168.875 116.615 169.685 ;
        RECT 115.385 168.705 116.615 168.875 ;
        RECT 116.785 169.305 117.170 170.275 ;
        RECT 117.340 169.985 117.665 170.445 ;
        RECT 118.185 169.815 118.465 170.275 ;
        RECT 117.340 169.595 118.465 169.815 ;
        RECT 115.365 167.895 115.875 168.430 ;
        RECT 116.095 168.100 116.340 168.705 ;
        RECT 116.785 168.635 117.065 169.305 ;
        RECT 117.340 169.135 117.790 169.595 ;
        RECT 118.655 169.425 119.055 170.275 ;
        RECT 119.455 169.985 119.725 170.445 ;
        RECT 119.895 169.815 120.180 170.275 ;
        RECT 117.235 168.805 117.790 169.135 ;
        RECT 117.960 168.865 119.055 169.425 ;
        RECT 117.340 168.695 117.790 168.805 ;
        RECT 116.785 168.065 117.170 168.635 ;
        RECT 117.340 168.525 118.465 168.695 ;
        RECT 117.340 167.895 117.665 168.355 ;
        RECT 118.185 168.065 118.465 168.525 ;
        RECT 118.655 168.065 119.055 168.865 ;
        RECT 119.225 169.595 120.180 169.815 ;
        RECT 119.225 168.695 119.435 169.595 ;
        RECT 120.555 169.515 120.725 170.275 ;
        RECT 120.905 169.685 121.235 170.445 ;
        RECT 119.605 168.865 120.295 169.425 ;
        RECT 120.555 169.345 121.220 169.515 ;
        RECT 121.405 169.370 121.675 170.275 ;
        RECT 121.850 170.020 122.185 170.445 ;
        RECT 122.355 169.840 122.540 170.245 ;
        RECT 121.050 169.200 121.220 169.345 ;
        RECT 120.485 168.795 120.815 169.165 ;
        RECT 121.050 168.870 121.335 169.200 ;
        RECT 119.225 168.525 120.180 168.695 ;
        RECT 121.050 168.615 121.220 168.870 ;
        RECT 119.455 167.895 119.725 168.355 ;
        RECT 119.895 168.065 120.180 168.525 ;
        RECT 120.555 168.445 121.220 168.615 ;
        RECT 121.505 168.570 121.675 169.370 ;
        RECT 120.555 168.065 120.725 168.445 ;
        RECT 120.905 167.895 121.235 168.275 ;
        RECT 121.415 168.065 121.675 168.570 ;
        RECT 121.875 169.665 122.540 169.840 ;
        RECT 122.745 169.665 123.075 170.445 ;
        RECT 121.875 168.635 122.215 169.665 ;
        RECT 123.245 169.475 123.515 170.245 ;
        RECT 122.385 169.305 123.515 169.475 ;
        RECT 122.385 168.805 122.635 169.305 ;
        RECT 121.875 168.465 122.560 168.635 ;
        RECT 122.815 168.555 123.175 169.135 ;
        RECT 121.850 167.895 122.185 168.295 ;
        RECT 122.355 168.065 122.560 168.465 ;
        RECT 123.345 168.395 123.515 169.305 ;
        RECT 123.685 169.355 126.275 170.445 ;
        RECT 126.445 169.355 127.655 170.445 ;
        RECT 123.685 168.835 124.895 169.355 ;
        RECT 125.065 168.665 126.275 169.185 ;
        RECT 126.445 168.815 126.965 169.355 ;
        RECT 122.770 167.895 123.045 168.375 ;
        RECT 123.255 168.065 123.515 168.395 ;
        RECT 123.685 167.895 126.275 168.665 ;
        RECT 127.135 168.645 127.655 169.185 ;
        RECT 126.445 167.895 127.655 168.645 ;
        RECT 14.580 167.725 127.740 167.895 ;
        RECT 14.665 166.975 15.875 167.725 ;
        RECT 14.665 166.435 15.185 166.975 ;
        RECT 16.045 166.955 17.715 167.725 ;
        RECT 17.890 167.180 23.235 167.725 ;
        RECT 15.355 166.265 15.875 166.805 ;
        RECT 14.665 165.175 15.875 166.265 ;
        RECT 16.045 166.265 16.795 166.785 ;
        RECT 16.965 166.435 17.715 166.955 ;
        RECT 16.045 165.175 17.715 166.265 ;
        RECT 19.480 165.610 19.830 166.860 ;
        RECT 21.310 166.350 21.650 167.180 ;
        RECT 23.410 167.175 23.665 167.465 ;
        RECT 23.835 167.345 24.165 167.725 ;
        RECT 23.410 167.005 24.160 167.175 ;
        RECT 23.410 166.185 23.760 166.835 ;
        RECT 23.930 166.015 24.160 167.005 ;
        RECT 23.410 165.845 24.160 166.015 ;
        RECT 17.890 165.175 23.235 165.610 ;
        RECT 23.410 165.345 23.665 165.845 ;
        RECT 23.835 165.175 24.165 165.675 ;
        RECT 24.335 165.345 24.505 167.465 ;
        RECT 24.865 167.365 25.195 167.725 ;
        RECT 25.365 167.335 25.860 167.505 ;
        RECT 26.065 167.335 26.920 167.505 ;
        RECT 24.735 166.145 25.195 167.195 ;
        RECT 24.675 165.360 25.000 166.145 ;
        RECT 25.365 165.975 25.535 167.335 ;
        RECT 25.705 166.425 26.055 167.045 ;
        RECT 26.225 166.825 26.580 167.045 ;
        RECT 26.225 166.235 26.395 166.825 ;
        RECT 26.750 166.625 26.920 167.335 ;
        RECT 27.795 167.265 28.125 167.725 ;
        RECT 28.335 167.365 28.685 167.535 ;
        RECT 27.125 166.795 27.915 167.045 ;
        RECT 28.335 166.975 28.595 167.365 ;
        RECT 28.905 167.275 29.855 167.555 ;
        RECT 30.025 167.285 30.215 167.725 ;
        RECT 30.385 167.345 31.455 167.515 ;
        RECT 28.085 166.625 28.255 166.805 ;
        RECT 25.365 165.805 25.760 165.975 ;
        RECT 25.930 165.845 26.395 166.235 ;
        RECT 26.565 166.455 28.255 166.625 ;
        RECT 25.590 165.675 25.760 165.805 ;
        RECT 26.565 165.675 26.735 166.455 ;
        RECT 28.425 166.285 28.595 166.975 ;
        RECT 27.095 166.115 28.595 166.285 ;
        RECT 28.785 166.315 28.995 167.105 ;
        RECT 29.165 166.485 29.515 167.105 ;
        RECT 29.685 166.495 29.855 167.275 ;
        RECT 30.385 167.115 30.555 167.345 ;
        RECT 30.025 166.945 30.555 167.115 ;
        RECT 30.025 166.665 30.245 166.945 ;
        RECT 30.725 166.775 30.965 167.175 ;
        RECT 29.685 166.325 30.090 166.495 ;
        RECT 30.425 166.405 30.965 166.775 ;
        RECT 31.135 166.990 31.455 167.345 ;
        RECT 31.700 167.265 32.005 167.725 ;
        RECT 32.175 167.015 32.430 167.545 ;
        RECT 31.135 166.815 31.460 166.990 ;
        RECT 31.135 166.515 32.050 166.815 ;
        RECT 31.310 166.485 32.050 166.515 ;
        RECT 28.785 166.155 29.460 166.315 ;
        RECT 29.920 166.235 30.090 166.325 ;
        RECT 28.785 166.145 29.750 166.155 ;
        RECT 28.425 165.975 28.595 166.115 ;
        RECT 25.170 165.175 25.420 165.635 ;
        RECT 25.590 165.345 25.840 165.675 ;
        RECT 26.055 165.345 26.735 165.675 ;
        RECT 26.905 165.775 27.980 165.945 ;
        RECT 28.425 165.805 28.985 165.975 ;
        RECT 29.290 165.855 29.750 166.145 ;
        RECT 29.920 166.065 31.140 166.235 ;
        RECT 26.905 165.435 27.075 165.775 ;
        RECT 27.310 165.175 27.640 165.605 ;
        RECT 27.810 165.435 27.980 165.775 ;
        RECT 28.275 165.175 28.645 165.635 ;
        RECT 28.815 165.345 28.985 165.805 ;
        RECT 29.920 165.685 30.090 166.065 ;
        RECT 31.310 165.895 31.480 166.485 ;
        RECT 32.220 166.365 32.430 167.015 ;
        RECT 29.220 165.345 30.090 165.685 ;
        RECT 30.680 165.725 31.480 165.895 ;
        RECT 30.260 165.175 30.510 165.635 ;
        RECT 30.680 165.435 30.850 165.725 ;
        RECT 31.030 165.175 31.360 165.555 ;
        RECT 31.700 165.175 32.005 166.315 ;
        RECT 32.175 165.485 32.430 166.365 ;
        RECT 32.605 167.050 32.865 167.555 ;
        RECT 33.045 167.345 33.375 167.725 ;
        RECT 33.555 167.175 33.725 167.555 ;
        RECT 34.085 167.260 34.335 167.725 ;
        RECT 32.605 166.250 32.775 167.050 ;
        RECT 33.060 167.005 33.725 167.175 ;
        RECT 34.505 167.085 34.675 167.555 ;
        RECT 34.925 167.265 35.095 167.725 ;
        RECT 35.345 167.085 35.515 167.555 ;
        RECT 35.765 167.265 35.935 167.725 ;
        RECT 36.185 167.085 36.355 167.555 ;
        RECT 36.725 167.265 36.990 167.725 ;
        RECT 33.060 166.750 33.230 167.005 ;
        RECT 33.985 166.905 36.355 167.085 ;
        RECT 37.205 167.000 37.495 167.725 ;
        RECT 37.705 166.905 37.935 167.725 ;
        RECT 38.105 166.925 38.435 167.555 ;
        RECT 32.945 166.420 33.230 166.750 ;
        RECT 33.465 166.455 33.795 166.825 ;
        RECT 33.060 166.275 33.230 166.420 ;
        RECT 33.985 166.315 34.335 166.905 ;
        RECT 34.505 166.485 37.015 166.735 ;
        RECT 37.685 166.485 38.015 166.735 ;
        RECT 32.605 165.345 32.875 166.250 ;
        RECT 33.060 166.105 33.725 166.275 ;
        RECT 33.985 166.145 36.435 166.315 ;
        RECT 33.985 166.125 34.755 166.145 ;
        RECT 33.045 165.175 33.375 165.935 ;
        RECT 33.555 165.345 33.725 166.105 ;
        RECT 34.085 165.175 34.255 165.635 ;
        RECT 34.425 165.345 34.755 166.125 ;
        RECT 34.925 165.175 35.095 165.975 ;
        RECT 35.265 165.345 35.595 166.145 ;
        RECT 35.765 165.175 35.935 165.975 ;
        RECT 36.105 165.345 36.435 166.145 ;
        RECT 36.695 165.175 36.990 166.315 ;
        RECT 37.205 165.175 37.495 166.340 ;
        RECT 38.185 166.325 38.435 166.925 ;
        RECT 38.605 166.905 38.815 167.725 ;
        RECT 39.160 167.095 39.445 167.555 ;
        RECT 39.615 167.265 39.885 167.725 ;
        RECT 39.160 166.925 40.115 167.095 ;
        RECT 37.705 165.175 37.935 166.315 ;
        RECT 38.105 165.345 38.435 166.325 ;
        RECT 38.605 165.175 38.815 166.315 ;
        RECT 39.045 166.195 39.735 166.755 ;
        RECT 39.905 166.025 40.115 166.925 ;
        RECT 39.160 165.805 40.115 166.025 ;
        RECT 40.285 166.755 40.685 167.555 ;
        RECT 40.875 167.095 41.155 167.555 ;
        RECT 41.675 167.265 42.000 167.725 ;
        RECT 40.875 166.925 42.000 167.095 ;
        RECT 42.170 166.985 42.555 167.555 ;
        RECT 41.550 166.815 42.000 166.925 ;
        RECT 40.285 166.195 41.380 166.755 ;
        RECT 41.550 166.485 42.105 166.815 ;
        RECT 39.160 165.345 39.445 165.805 ;
        RECT 39.615 165.175 39.885 165.635 ;
        RECT 40.285 165.345 40.685 166.195 ;
        RECT 41.550 166.025 42.000 166.485 ;
        RECT 42.275 166.315 42.555 166.985 ;
        RECT 40.875 165.805 42.000 166.025 ;
        RECT 40.875 165.345 41.155 165.805 ;
        RECT 41.675 165.175 42.000 165.635 ;
        RECT 42.170 165.345 42.555 166.315 ;
        RECT 42.725 166.985 43.110 167.555 ;
        RECT 43.280 167.265 43.605 167.725 ;
        RECT 44.125 167.095 44.405 167.555 ;
        RECT 42.725 166.315 43.005 166.985 ;
        RECT 43.280 166.925 44.405 167.095 ;
        RECT 43.280 166.815 43.730 166.925 ;
        RECT 43.175 166.485 43.730 166.815 ;
        RECT 44.595 166.755 44.995 167.555 ;
        RECT 45.395 167.265 45.665 167.725 ;
        RECT 45.835 167.095 46.120 167.555 ;
        RECT 42.725 165.345 43.110 166.315 ;
        RECT 43.280 166.025 43.730 166.485 ;
        RECT 43.900 166.195 44.995 166.755 ;
        RECT 43.280 165.805 44.405 166.025 ;
        RECT 43.280 165.175 43.605 165.635 ;
        RECT 44.125 165.345 44.405 165.805 ;
        RECT 44.595 165.345 44.995 166.195 ;
        RECT 45.165 166.925 46.120 167.095 ;
        RECT 47.330 167.015 47.585 167.545 ;
        RECT 47.755 167.265 48.060 167.725 ;
        RECT 48.305 167.345 49.375 167.515 ;
        RECT 45.165 166.025 45.375 166.925 ;
        RECT 45.545 166.195 46.235 166.755 ;
        RECT 47.330 166.365 47.540 167.015 ;
        RECT 48.305 166.990 48.625 167.345 ;
        RECT 48.300 166.815 48.625 166.990 ;
        RECT 47.710 166.515 48.625 166.815 ;
        RECT 48.795 166.775 49.035 167.175 ;
        RECT 49.205 167.115 49.375 167.345 ;
        RECT 49.545 167.285 49.735 167.725 ;
        RECT 49.905 167.275 50.855 167.555 ;
        RECT 51.075 167.365 51.425 167.535 ;
        RECT 49.205 166.945 49.735 167.115 ;
        RECT 47.710 166.485 48.450 166.515 ;
        RECT 45.165 165.805 46.120 166.025 ;
        RECT 45.395 165.175 45.665 165.635 ;
        RECT 45.835 165.345 46.120 165.805 ;
        RECT 47.330 165.485 47.585 166.365 ;
        RECT 47.755 165.175 48.060 166.315 ;
        RECT 48.280 165.895 48.450 166.485 ;
        RECT 48.795 166.405 49.335 166.775 ;
        RECT 49.515 166.665 49.735 166.945 ;
        RECT 49.905 166.495 50.075 167.275 ;
        RECT 49.670 166.325 50.075 166.495 ;
        RECT 50.245 166.485 50.595 167.105 ;
        RECT 49.670 166.235 49.840 166.325 ;
        RECT 50.765 166.315 50.975 167.105 ;
        RECT 48.620 166.065 49.840 166.235 ;
        RECT 50.300 166.155 50.975 166.315 ;
        RECT 48.280 165.725 49.080 165.895 ;
        RECT 48.400 165.175 48.730 165.555 ;
        RECT 48.910 165.435 49.080 165.725 ;
        RECT 49.670 165.685 49.840 166.065 ;
        RECT 50.010 166.145 50.975 166.155 ;
        RECT 51.165 166.975 51.425 167.365 ;
        RECT 51.635 167.265 51.965 167.725 ;
        RECT 52.840 167.335 53.695 167.505 ;
        RECT 53.900 167.335 54.395 167.505 ;
        RECT 54.565 167.365 54.895 167.725 ;
        RECT 51.165 166.285 51.335 166.975 ;
        RECT 51.505 166.625 51.675 166.805 ;
        RECT 51.845 166.795 52.635 167.045 ;
        RECT 52.840 166.625 53.010 167.335 ;
        RECT 53.180 166.825 53.535 167.045 ;
        RECT 51.505 166.455 53.195 166.625 ;
        RECT 50.010 165.855 50.470 166.145 ;
        RECT 51.165 166.115 52.665 166.285 ;
        RECT 51.165 165.975 51.335 166.115 ;
        RECT 50.775 165.805 51.335 165.975 ;
        RECT 49.250 165.175 49.500 165.635 ;
        RECT 49.670 165.345 50.540 165.685 ;
        RECT 50.775 165.345 50.945 165.805 ;
        RECT 51.780 165.775 52.855 165.945 ;
        RECT 51.115 165.175 51.485 165.635 ;
        RECT 51.780 165.435 51.950 165.775 ;
        RECT 52.120 165.175 52.450 165.605 ;
        RECT 52.685 165.435 52.855 165.775 ;
        RECT 53.025 165.675 53.195 166.455 ;
        RECT 53.365 166.235 53.535 166.825 ;
        RECT 53.705 166.425 54.055 167.045 ;
        RECT 53.365 165.845 53.830 166.235 ;
        RECT 54.225 165.975 54.395 167.335 ;
        RECT 54.565 166.145 55.025 167.195 ;
        RECT 54.000 165.805 54.395 165.975 ;
        RECT 54.000 165.675 54.170 165.805 ;
        RECT 53.025 165.345 53.705 165.675 ;
        RECT 53.920 165.345 54.170 165.675 ;
        RECT 54.340 165.175 54.590 165.635 ;
        RECT 54.760 165.360 55.085 166.145 ;
        RECT 55.255 165.345 55.425 167.465 ;
        RECT 55.595 167.345 55.925 167.725 ;
        RECT 56.095 167.175 56.350 167.465 ;
        RECT 55.600 167.005 56.350 167.175 ;
        RECT 55.600 166.015 55.830 167.005 ;
        RECT 56.525 166.955 58.195 167.725 ;
        RECT 56.000 166.185 56.350 166.835 ;
        RECT 56.525 166.265 57.275 166.785 ;
        RECT 57.445 166.435 58.195 166.955 ;
        RECT 58.425 166.905 58.635 167.725 ;
        RECT 58.805 166.925 59.135 167.555 ;
        RECT 58.805 166.325 59.055 166.925 ;
        RECT 59.305 166.905 59.535 167.725 ;
        RECT 60.355 166.925 60.685 167.725 ;
        RECT 60.855 167.075 61.025 167.555 ;
        RECT 61.195 167.245 61.525 167.725 ;
        RECT 61.695 167.075 61.865 167.555 ;
        RECT 62.115 167.245 62.355 167.725 ;
        RECT 62.535 167.075 62.705 167.555 ;
        RECT 60.855 166.905 61.865 167.075 ;
        RECT 62.070 166.905 62.705 167.075 ;
        RECT 62.965 167.000 63.255 167.725 ;
        RECT 63.425 166.955 65.095 167.725 ;
        RECT 65.325 167.245 65.605 167.725 ;
        RECT 65.775 167.075 66.035 167.465 ;
        RECT 66.210 167.245 66.465 167.725 ;
        RECT 66.635 167.075 66.930 167.465 ;
        RECT 67.110 167.245 67.385 167.725 ;
        RECT 67.555 167.225 67.855 167.555 ;
        RECT 59.225 166.485 59.555 166.735 ;
        RECT 60.855 166.705 61.350 166.905 ;
        RECT 62.070 166.735 62.240 166.905 ;
        RECT 60.855 166.535 61.355 166.705 ;
        RECT 61.740 166.565 62.240 166.735 ;
        RECT 60.855 166.365 61.350 166.535 ;
        RECT 55.600 165.845 56.350 166.015 ;
        RECT 55.595 165.175 55.925 165.675 ;
        RECT 56.095 165.345 56.350 165.845 ;
        RECT 56.525 165.175 58.195 166.265 ;
        RECT 58.425 165.175 58.635 166.315 ;
        RECT 58.805 165.345 59.135 166.325 ;
        RECT 59.305 165.175 59.535 166.315 ;
        RECT 60.355 165.175 60.685 166.325 ;
        RECT 60.855 166.195 61.865 166.365 ;
        RECT 60.855 165.345 61.025 166.195 ;
        RECT 61.195 165.175 61.525 165.975 ;
        RECT 61.695 165.345 61.865 166.195 ;
        RECT 62.070 166.325 62.240 166.565 ;
        RECT 62.410 166.495 62.790 166.735 ;
        RECT 62.070 166.155 62.785 166.325 ;
        RECT 62.045 165.175 62.285 165.975 ;
        RECT 62.455 165.345 62.785 166.155 ;
        RECT 62.965 165.175 63.255 166.340 ;
        RECT 63.425 166.265 64.175 166.785 ;
        RECT 64.345 166.435 65.095 166.955 ;
        RECT 65.280 166.905 66.930 167.075 ;
        RECT 65.280 166.395 65.685 166.905 ;
        RECT 65.855 166.565 66.995 166.735 ;
        RECT 63.425 165.175 65.095 166.265 ;
        RECT 65.280 166.225 66.035 166.395 ;
        RECT 65.320 165.175 65.605 166.045 ;
        RECT 65.775 165.975 66.035 166.225 ;
        RECT 66.825 166.315 66.995 166.565 ;
        RECT 67.165 166.485 67.515 167.055 ;
        RECT 67.685 166.315 67.855 167.225 ;
        RECT 66.825 166.145 67.855 166.315 ;
        RECT 65.775 165.805 66.895 165.975 ;
        RECT 65.775 165.345 66.035 165.805 ;
        RECT 66.210 165.175 66.465 165.635 ;
        RECT 66.635 165.345 66.895 165.805 ;
        RECT 67.065 165.175 67.375 165.975 ;
        RECT 67.545 165.345 67.855 166.145 ;
        RECT 68.025 167.225 68.325 167.555 ;
        RECT 68.495 167.245 68.770 167.725 ;
        RECT 68.025 166.315 68.195 167.225 ;
        RECT 68.950 167.075 69.245 167.465 ;
        RECT 69.415 167.245 69.670 167.725 ;
        RECT 69.845 167.075 70.105 167.465 ;
        RECT 70.275 167.245 70.555 167.725 ;
        RECT 70.795 167.195 71.125 167.555 ;
        RECT 71.295 167.365 71.625 167.725 ;
        RECT 71.825 167.195 72.155 167.555 ;
        RECT 68.365 166.485 68.715 167.055 ;
        RECT 68.950 166.905 70.600 167.075 ;
        RECT 70.795 166.985 72.155 167.195 ;
        RECT 72.665 166.965 73.375 167.555 ;
        RECT 68.885 166.565 70.025 166.735 ;
        RECT 68.885 166.315 69.055 166.565 ;
        RECT 70.195 166.395 70.600 166.905 ;
        RECT 73.145 166.875 73.375 166.965 ;
        RECT 73.545 166.955 75.215 167.725 ;
        RECT 70.785 166.485 71.095 166.815 ;
        RECT 71.305 166.485 71.680 166.815 ;
        RECT 72.000 166.485 72.495 166.815 ;
        RECT 68.025 166.145 69.055 166.315 ;
        RECT 69.845 166.225 70.600 166.395 ;
        RECT 68.025 165.345 68.335 166.145 ;
        RECT 69.845 165.975 70.105 166.225 ;
        RECT 68.505 165.175 68.815 165.975 ;
        RECT 68.985 165.805 70.105 165.975 ;
        RECT 68.985 165.345 69.245 165.805 ;
        RECT 69.415 165.175 69.670 165.635 ;
        RECT 69.845 165.345 70.105 165.805 ;
        RECT 70.275 165.175 70.560 166.045 ;
        RECT 70.795 165.175 71.125 166.235 ;
        RECT 71.305 165.560 71.475 166.485 ;
        RECT 71.645 165.995 71.975 166.215 ;
        RECT 72.170 166.195 72.495 166.485 ;
        RECT 72.670 166.195 73.000 166.735 ;
        RECT 73.170 165.995 73.375 166.875 ;
        RECT 71.645 165.765 73.375 165.995 ;
        RECT 71.645 165.365 71.975 165.765 ;
        RECT 72.145 165.175 72.475 165.535 ;
        RECT 72.675 165.345 73.375 165.765 ;
        RECT 73.545 166.265 74.295 166.785 ;
        RECT 74.465 166.435 75.215 166.955 ;
        RECT 75.760 167.015 76.015 167.545 ;
        RECT 76.195 167.265 76.480 167.725 ;
        RECT 73.545 165.175 75.215 166.265 ;
        RECT 75.760 166.155 75.940 167.015 ;
        RECT 76.660 166.815 76.910 167.465 ;
        RECT 76.110 166.485 76.910 166.815 ;
        RECT 75.760 165.685 76.015 166.155 ;
        RECT 75.675 165.515 76.015 165.685 ;
        RECT 75.760 165.485 76.015 165.515 ;
        RECT 76.195 165.175 76.480 165.975 ;
        RECT 76.660 165.895 76.910 166.485 ;
        RECT 77.110 167.130 77.430 167.460 ;
        RECT 77.610 167.245 78.270 167.725 ;
        RECT 78.470 167.335 79.320 167.505 ;
        RECT 77.110 166.235 77.300 167.130 ;
        RECT 77.620 166.805 78.280 167.075 ;
        RECT 77.950 166.745 78.280 166.805 ;
        RECT 77.470 166.575 77.800 166.635 ;
        RECT 78.470 166.575 78.640 167.335 ;
        RECT 79.880 167.265 80.200 167.725 ;
        RECT 80.400 167.085 80.650 167.515 ;
        RECT 80.940 167.285 81.350 167.725 ;
        RECT 81.520 167.345 82.535 167.545 ;
        RECT 78.810 166.915 80.060 167.085 ;
        RECT 78.810 166.795 79.140 166.915 ;
        RECT 77.470 166.405 79.370 166.575 ;
        RECT 77.110 166.065 79.030 166.235 ;
        RECT 77.110 166.045 77.430 166.065 ;
        RECT 76.660 165.385 76.990 165.895 ;
        RECT 77.260 165.435 77.430 166.045 ;
        RECT 79.200 165.895 79.370 166.405 ;
        RECT 79.540 166.335 79.720 166.745 ;
        RECT 79.890 166.155 80.060 166.915 ;
        RECT 77.600 165.175 77.930 165.865 ;
        RECT 78.160 165.725 79.370 165.895 ;
        RECT 79.540 165.845 80.060 166.155 ;
        RECT 80.230 166.745 80.650 167.085 ;
        RECT 80.940 166.745 81.350 167.075 ;
        RECT 80.230 165.975 80.420 166.745 ;
        RECT 81.520 166.615 81.690 167.345 ;
        RECT 82.835 167.175 83.005 167.505 ;
        RECT 83.175 167.345 83.505 167.725 ;
        RECT 81.860 166.795 82.210 167.165 ;
        RECT 81.520 166.575 81.940 166.615 ;
        RECT 80.590 166.405 81.940 166.575 ;
        RECT 80.590 166.245 80.840 166.405 ;
        RECT 81.350 165.975 81.600 166.235 ;
        RECT 80.230 165.725 81.600 165.975 ;
        RECT 78.160 165.435 78.400 165.725 ;
        RECT 79.200 165.645 79.370 165.725 ;
        RECT 78.600 165.175 79.020 165.555 ;
        RECT 79.200 165.395 79.830 165.645 ;
        RECT 80.300 165.175 80.630 165.555 ;
        RECT 80.800 165.435 80.970 165.725 ;
        RECT 81.770 165.560 81.940 166.405 ;
        RECT 82.390 166.235 82.610 167.105 ;
        RECT 82.835 166.985 83.530 167.175 ;
        RECT 82.110 165.855 82.610 166.235 ;
        RECT 82.780 166.185 83.190 166.805 ;
        RECT 83.360 166.015 83.530 166.985 ;
        RECT 82.835 165.845 83.530 166.015 ;
        RECT 81.150 165.175 81.530 165.555 ;
        RECT 81.770 165.390 82.600 165.560 ;
        RECT 82.835 165.345 83.005 165.845 ;
        RECT 83.175 165.175 83.505 165.675 ;
        RECT 83.720 165.345 83.945 167.465 ;
        RECT 84.115 167.345 84.445 167.725 ;
        RECT 84.615 167.175 84.785 167.465 ;
        RECT 84.120 167.005 84.785 167.175 ;
        RECT 84.120 166.015 84.350 167.005 ;
        RECT 85.105 166.905 85.315 167.725 ;
        RECT 85.485 166.925 85.815 167.555 ;
        RECT 84.520 166.185 84.870 166.835 ;
        RECT 85.485 166.325 85.735 166.925 ;
        RECT 85.985 166.905 86.215 167.725 ;
        RECT 86.485 166.905 86.695 167.725 ;
        RECT 86.865 166.925 87.195 167.555 ;
        RECT 85.905 166.485 86.235 166.735 ;
        RECT 86.865 166.325 87.115 166.925 ;
        RECT 87.365 166.905 87.595 167.725 ;
        RECT 88.725 167.000 89.015 167.725 ;
        RECT 89.645 166.955 93.155 167.725 ;
        RECT 87.285 166.485 87.615 166.735 ;
        RECT 84.120 165.845 84.785 166.015 ;
        RECT 84.115 165.175 84.445 165.675 ;
        RECT 84.615 165.345 84.785 165.845 ;
        RECT 85.105 165.175 85.315 166.315 ;
        RECT 85.485 165.345 85.815 166.325 ;
        RECT 85.985 165.175 86.215 166.315 ;
        RECT 86.485 165.175 86.695 166.315 ;
        RECT 86.865 165.345 87.195 166.325 ;
        RECT 87.365 165.175 87.595 166.315 ;
        RECT 88.725 165.175 89.015 166.340 ;
        RECT 89.645 166.265 91.335 166.785 ;
        RECT 91.505 166.435 93.155 166.955 ;
        RECT 93.600 166.915 93.845 167.520 ;
        RECT 94.065 167.190 94.575 167.725 ;
        RECT 93.325 166.745 94.555 166.915 ;
        RECT 89.645 165.175 93.155 166.265 ;
        RECT 93.325 165.935 93.665 166.745 ;
        RECT 93.835 166.180 94.585 166.370 ;
        RECT 93.325 165.525 93.840 165.935 ;
        RECT 94.075 165.175 94.245 165.935 ;
        RECT 94.415 165.515 94.585 166.180 ;
        RECT 94.755 166.195 94.945 167.555 ;
        RECT 95.115 166.705 95.390 167.555 ;
        RECT 95.580 167.190 96.110 167.555 ;
        RECT 96.535 167.325 96.865 167.725 ;
        RECT 95.935 167.155 96.110 167.190 ;
        RECT 95.115 166.535 95.395 166.705 ;
        RECT 95.115 166.395 95.390 166.535 ;
        RECT 95.595 166.195 95.765 166.995 ;
        RECT 94.755 166.025 95.765 166.195 ;
        RECT 95.935 166.985 96.865 167.155 ;
        RECT 97.035 166.985 97.290 167.555 ;
        RECT 95.935 165.855 96.105 166.985 ;
        RECT 96.695 166.815 96.865 166.985 ;
        RECT 94.980 165.685 96.105 165.855 ;
        RECT 96.275 166.485 96.470 166.815 ;
        RECT 96.695 166.485 96.950 166.815 ;
        RECT 96.275 165.515 96.445 166.485 ;
        RECT 97.120 166.315 97.290 166.985 ;
        RECT 97.840 167.015 98.095 167.545 ;
        RECT 98.275 167.265 98.560 167.725 ;
        RECT 97.840 166.365 98.020 167.015 ;
        RECT 98.740 166.815 98.990 167.465 ;
        RECT 98.190 166.485 98.990 166.815 ;
        RECT 94.415 165.345 96.445 165.515 ;
        RECT 96.615 165.175 96.785 166.315 ;
        RECT 96.955 165.345 97.290 166.315 ;
        RECT 97.755 166.195 98.020 166.365 ;
        RECT 97.840 166.155 98.020 166.195 ;
        RECT 97.840 165.485 98.095 166.155 ;
        RECT 98.275 165.175 98.560 165.975 ;
        RECT 98.740 165.895 98.990 166.485 ;
        RECT 99.190 167.130 99.510 167.460 ;
        RECT 99.690 167.245 100.350 167.725 ;
        RECT 100.550 167.335 101.400 167.505 ;
        RECT 99.190 166.235 99.380 167.130 ;
        RECT 99.700 166.805 100.360 167.075 ;
        RECT 100.030 166.745 100.360 166.805 ;
        RECT 99.550 166.575 99.880 166.635 ;
        RECT 100.550 166.575 100.720 167.335 ;
        RECT 101.960 167.265 102.280 167.725 ;
        RECT 102.480 167.085 102.730 167.515 ;
        RECT 103.020 167.285 103.430 167.725 ;
        RECT 103.600 167.345 104.615 167.545 ;
        RECT 100.890 166.915 102.140 167.085 ;
        RECT 100.890 166.795 101.220 166.915 ;
        RECT 99.550 166.405 101.450 166.575 ;
        RECT 99.190 166.065 101.110 166.235 ;
        RECT 99.190 166.045 99.510 166.065 ;
        RECT 98.740 165.385 99.070 165.895 ;
        RECT 99.340 165.435 99.510 166.045 ;
        RECT 101.280 165.895 101.450 166.405 ;
        RECT 101.620 166.335 101.800 166.745 ;
        RECT 101.970 166.155 102.140 166.915 ;
        RECT 99.680 165.175 100.010 165.865 ;
        RECT 100.240 165.725 101.450 165.895 ;
        RECT 101.620 165.845 102.140 166.155 ;
        RECT 102.310 166.745 102.730 167.085 ;
        RECT 103.020 166.745 103.430 167.075 ;
        RECT 102.310 165.975 102.500 166.745 ;
        RECT 103.600 166.615 103.770 167.345 ;
        RECT 104.915 167.175 105.085 167.505 ;
        RECT 105.255 167.345 105.585 167.725 ;
        RECT 103.940 166.795 104.290 167.165 ;
        RECT 103.600 166.575 104.020 166.615 ;
        RECT 102.670 166.405 104.020 166.575 ;
        RECT 102.670 166.245 102.920 166.405 ;
        RECT 103.430 165.975 103.680 166.235 ;
        RECT 102.310 165.725 103.680 165.975 ;
        RECT 100.240 165.435 100.480 165.725 ;
        RECT 101.280 165.645 101.450 165.725 ;
        RECT 100.680 165.175 101.100 165.555 ;
        RECT 101.280 165.395 101.910 165.645 ;
        RECT 102.380 165.175 102.710 165.555 ;
        RECT 102.880 165.435 103.050 165.725 ;
        RECT 103.850 165.560 104.020 166.405 ;
        RECT 104.470 166.235 104.690 167.105 ;
        RECT 104.915 166.985 105.610 167.175 ;
        RECT 104.190 165.855 104.690 166.235 ;
        RECT 104.860 166.185 105.270 166.805 ;
        RECT 105.440 166.015 105.610 166.985 ;
        RECT 104.915 165.845 105.610 166.015 ;
        RECT 103.230 165.175 103.610 165.555 ;
        RECT 103.850 165.390 104.680 165.560 ;
        RECT 104.915 165.345 105.085 165.845 ;
        RECT 105.255 165.175 105.585 165.675 ;
        RECT 105.800 165.345 106.025 167.465 ;
        RECT 106.195 167.345 106.525 167.725 ;
        RECT 106.695 167.175 106.865 167.465 ;
        RECT 106.200 167.005 106.865 167.175 ;
        RECT 107.240 167.095 107.525 167.555 ;
        RECT 107.695 167.265 107.965 167.725 ;
        RECT 106.200 166.015 106.430 167.005 ;
        RECT 107.240 166.925 108.195 167.095 ;
        RECT 106.600 166.185 106.950 166.835 ;
        RECT 107.125 166.195 107.815 166.755 ;
        RECT 107.985 166.025 108.195 166.925 ;
        RECT 106.200 165.845 106.865 166.015 ;
        RECT 106.195 165.175 106.525 165.675 ;
        RECT 106.695 165.345 106.865 165.845 ;
        RECT 107.240 165.805 108.195 166.025 ;
        RECT 108.365 166.755 108.765 167.555 ;
        RECT 108.955 167.095 109.235 167.555 ;
        RECT 109.755 167.265 110.080 167.725 ;
        RECT 108.955 166.925 110.080 167.095 ;
        RECT 110.250 166.985 110.635 167.555 ;
        RECT 109.630 166.815 110.080 166.925 ;
        RECT 108.365 166.195 109.460 166.755 ;
        RECT 109.630 166.485 110.185 166.815 ;
        RECT 107.240 165.345 107.525 165.805 ;
        RECT 107.695 165.175 107.965 165.635 ;
        RECT 108.365 165.345 108.765 166.195 ;
        RECT 109.630 166.025 110.080 166.485 ;
        RECT 110.355 166.315 110.635 166.985 ;
        RECT 110.920 167.095 111.205 167.555 ;
        RECT 111.375 167.265 111.645 167.725 ;
        RECT 110.920 166.925 111.875 167.095 ;
        RECT 108.955 165.805 110.080 166.025 ;
        RECT 108.955 165.345 109.235 165.805 ;
        RECT 109.755 165.175 110.080 165.635 ;
        RECT 110.250 165.345 110.635 166.315 ;
        RECT 110.805 166.195 111.495 166.755 ;
        RECT 111.665 166.025 111.875 166.925 ;
        RECT 110.920 165.805 111.875 166.025 ;
        RECT 112.045 166.755 112.445 167.555 ;
        RECT 112.635 167.095 112.915 167.555 ;
        RECT 113.435 167.265 113.760 167.725 ;
        RECT 112.635 166.925 113.760 167.095 ;
        RECT 113.930 166.985 114.315 167.555 ;
        RECT 114.485 167.000 114.775 167.725 ;
        RECT 115.870 167.015 116.125 167.545 ;
        RECT 116.295 167.265 116.600 167.725 ;
        RECT 116.845 167.345 117.915 167.515 ;
        RECT 113.310 166.815 113.760 166.925 ;
        RECT 112.045 166.195 113.140 166.755 ;
        RECT 113.310 166.485 113.865 166.815 ;
        RECT 110.920 165.345 111.205 165.805 ;
        RECT 111.375 165.175 111.645 165.635 ;
        RECT 112.045 165.345 112.445 166.195 ;
        RECT 113.310 166.025 113.760 166.485 ;
        RECT 114.035 166.315 114.315 166.985 ;
        RECT 115.870 166.365 116.080 167.015 ;
        RECT 116.845 166.990 117.165 167.345 ;
        RECT 116.840 166.815 117.165 166.990 ;
        RECT 116.250 166.515 117.165 166.815 ;
        RECT 117.335 166.775 117.575 167.175 ;
        RECT 117.745 167.115 117.915 167.345 ;
        RECT 118.085 167.285 118.275 167.725 ;
        RECT 118.445 167.275 119.395 167.555 ;
        RECT 119.615 167.365 119.965 167.535 ;
        RECT 117.745 166.945 118.275 167.115 ;
        RECT 116.250 166.485 116.990 166.515 ;
        RECT 112.635 165.805 113.760 166.025 ;
        RECT 112.635 165.345 112.915 165.805 ;
        RECT 113.435 165.175 113.760 165.635 ;
        RECT 113.930 165.345 114.315 166.315 ;
        RECT 114.485 165.175 114.775 166.340 ;
        RECT 115.870 165.485 116.125 166.365 ;
        RECT 116.295 165.175 116.600 166.315 ;
        RECT 116.820 165.895 116.990 166.485 ;
        RECT 117.335 166.405 117.875 166.775 ;
        RECT 118.055 166.665 118.275 166.945 ;
        RECT 118.445 166.495 118.615 167.275 ;
        RECT 118.210 166.325 118.615 166.495 ;
        RECT 118.785 166.485 119.135 167.105 ;
        RECT 118.210 166.235 118.380 166.325 ;
        RECT 119.305 166.315 119.515 167.105 ;
        RECT 117.160 166.065 118.380 166.235 ;
        RECT 118.840 166.155 119.515 166.315 ;
        RECT 116.820 165.725 117.620 165.895 ;
        RECT 116.940 165.175 117.270 165.555 ;
        RECT 117.450 165.435 117.620 165.725 ;
        RECT 118.210 165.685 118.380 166.065 ;
        RECT 118.550 166.145 119.515 166.155 ;
        RECT 119.705 166.975 119.965 167.365 ;
        RECT 120.175 167.265 120.505 167.725 ;
        RECT 121.380 167.335 122.235 167.505 ;
        RECT 122.440 167.335 122.935 167.505 ;
        RECT 123.105 167.365 123.435 167.725 ;
        RECT 119.705 166.285 119.875 166.975 ;
        RECT 120.045 166.625 120.215 166.805 ;
        RECT 120.385 166.795 121.175 167.045 ;
        RECT 121.380 166.625 121.550 167.335 ;
        RECT 121.720 166.825 122.075 167.045 ;
        RECT 120.045 166.455 121.735 166.625 ;
        RECT 118.550 165.855 119.010 166.145 ;
        RECT 119.705 166.115 121.205 166.285 ;
        RECT 119.705 165.975 119.875 166.115 ;
        RECT 119.315 165.805 119.875 165.975 ;
        RECT 117.790 165.175 118.040 165.635 ;
        RECT 118.210 165.345 119.080 165.685 ;
        RECT 119.315 165.345 119.485 165.805 ;
        RECT 120.320 165.775 121.395 165.945 ;
        RECT 119.655 165.175 120.025 165.635 ;
        RECT 120.320 165.435 120.490 165.775 ;
        RECT 120.660 165.175 120.990 165.605 ;
        RECT 121.225 165.435 121.395 165.775 ;
        RECT 121.565 165.675 121.735 166.455 ;
        RECT 121.905 166.235 122.075 166.825 ;
        RECT 122.245 166.425 122.595 167.045 ;
        RECT 121.905 165.845 122.370 166.235 ;
        RECT 122.765 165.975 122.935 167.335 ;
        RECT 123.105 166.145 123.565 167.195 ;
        RECT 122.540 165.805 122.935 165.975 ;
        RECT 122.540 165.675 122.710 165.805 ;
        RECT 121.565 165.345 122.245 165.675 ;
        RECT 122.460 165.345 122.710 165.675 ;
        RECT 122.880 165.175 123.130 165.635 ;
        RECT 123.300 165.360 123.625 166.145 ;
        RECT 123.795 165.345 123.965 167.465 ;
        RECT 124.135 167.345 124.465 167.725 ;
        RECT 124.635 167.175 124.890 167.465 ;
        RECT 124.140 167.005 124.890 167.175 ;
        RECT 124.140 166.015 124.370 167.005 ;
        RECT 125.065 166.975 126.275 167.725 ;
        RECT 126.445 166.975 127.655 167.725 ;
        RECT 124.540 166.185 124.890 166.835 ;
        RECT 125.065 166.265 125.585 166.805 ;
        RECT 125.755 166.435 126.275 166.975 ;
        RECT 126.445 166.265 126.965 166.805 ;
        RECT 127.135 166.435 127.655 166.975 ;
        RECT 124.140 165.845 124.890 166.015 ;
        RECT 124.135 165.175 124.465 165.675 ;
        RECT 124.635 165.345 124.890 165.845 ;
        RECT 125.065 165.175 126.275 166.265 ;
        RECT 126.445 165.175 127.655 166.265 ;
        RECT 14.580 165.005 127.740 165.175 ;
        RECT 14.665 163.915 15.875 165.005 ;
        RECT 14.665 163.205 15.185 163.745 ;
        RECT 15.355 163.375 15.875 163.915 ;
        RECT 16.045 163.915 18.635 165.005 ;
        RECT 18.810 164.570 24.155 165.005 ;
        RECT 16.045 163.395 17.255 163.915 ;
        RECT 17.425 163.225 18.635 163.745 ;
        RECT 20.400 163.320 20.750 164.570 ;
        RECT 24.325 163.840 24.615 165.005 ;
        RECT 25.705 163.930 25.975 164.835 ;
        RECT 26.145 164.245 26.475 165.005 ;
        RECT 26.655 164.075 26.825 164.835 ;
        RECT 27.090 164.335 27.345 164.835 ;
        RECT 27.515 164.505 27.845 165.005 ;
        RECT 27.090 164.165 27.840 164.335 ;
        RECT 14.665 162.455 15.875 163.205 ;
        RECT 16.045 162.455 18.635 163.225 ;
        RECT 22.230 163.000 22.570 163.830 ;
        RECT 18.810 162.455 24.155 163.000 ;
        RECT 24.325 162.455 24.615 163.180 ;
        RECT 25.705 163.130 25.875 163.930 ;
        RECT 26.160 163.905 26.825 164.075 ;
        RECT 26.160 163.760 26.330 163.905 ;
        RECT 26.045 163.430 26.330 163.760 ;
        RECT 26.160 163.175 26.330 163.430 ;
        RECT 26.565 163.355 26.895 163.725 ;
        RECT 27.090 163.345 27.440 163.995 ;
        RECT 27.610 163.175 27.840 164.165 ;
        RECT 25.705 162.625 25.965 163.130 ;
        RECT 26.160 163.005 26.825 163.175 ;
        RECT 26.145 162.455 26.475 162.835 ;
        RECT 26.655 162.625 26.825 163.005 ;
        RECT 27.090 163.005 27.840 163.175 ;
        RECT 27.090 162.715 27.345 163.005 ;
        RECT 27.515 162.455 27.845 162.835 ;
        RECT 28.015 162.715 28.185 164.835 ;
        RECT 28.355 164.035 28.680 164.820 ;
        RECT 28.850 164.545 29.100 165.005 ;
        RECT 29.270 164.505 29.520 164.835 ;
        RECT 29.735 164.505 30.415 164.835 ;
        RECT 29.270 164.375 29.440 164.505 ;
        RECT 29.045 164.205 29.440 164.375 ;
        RECT 28.415 162.985 28.875 164.035 ;
        RECT 29.045 162.845 29.215 164.205 ;
        RECT 29.610 163.945 30.075 164.335 ;
        RECT 29.385 163.135 29.735 163.755 ;
        RECT 29.905 163.355 30.075 163.945 ;
        RECT 30.245 163.725 30.415 164.505 ;
        RECT 30.585 164.405 30.755 164.745 ;
        RECT 30.990 164.575 31.320 165.005 ;
        RECT 31.490 164.405 31.660 164.745 ;
        RECT 31.955 164.545 32.325 165.005 ;
        RECT 30.585 164.235 31.660 164.405 ;
        RECT 32.495 164.375 32.665 164.835 ;
        RECT 32.900 164.495 33.770 164.835 ;
        RECT 33.940 164.545 34.190 165.005 ;
        RECT 32.105 164.205 32.665 164.375 ;
        RECT 32.105 164.065 32.275 164.205 ;
        RECT 30.775 163.895 32.275 164.065 ;
        RECT 32.970 164.035 33.430 164.325 ;
        RECT 30.245 163.555 31.935 163.725 ;
        RECT 29.905 163.135 30.260 163.355 ;
        RECT 30.430 162.845 30.600 163.555 ;
        RECT 30.805 163.135 31.595 163.385 ;
        RECT 31.765 163.375 31.935 163.555 ;
        RECT 32.105 163.205 32.275 163.895 ;
        RECT 28.545 162.455 28.875 162.815 ;
        RECT 29.045 162.675 29.540 162.845 ;
        RECT 29.745 162.675 30.600 162.845 ;
        RECT 31.475 162.455 31.805 162.915 ;
        RECT 32.015 162.815 32.275 163.205 ;
        RECT 32.465 164.025 33.430 164.035 ;
        RECT 33.600 164.115 33.770 164.495 ;
        RECT 34.360 164.455 34.530 164.745 ;
        RECT 34.710 164.625 35.040 165.005 ;
        RECT 34.360 164.285 35.160 164.455 ;
        RECT 32.465 163.865 33.140 164.025 ;
        RECT 33.600 163.945 34.820 164.115 ;
        RECT 32.465 163.075 32.675 163.865 ;
        RECT 33.600 163.855 33.770 163.945 ;
        RECT 32.845 163.075 33.195 163.695 ;
        RECT 33.365 163.685 33.770 163.855 ;
        RECT 33.365 162.905 33.535 163.685 ;
        RECT 33.705 163.235 33.925 163.515 ;
        RECT 34.105 163.405 34.645 163.775 ;
        RECT 34.990 163.695 35.160 164.285 ;
        RECT 35.380 163.865 35.685 165.005 ;
        RECT 35.855 163.815 36.110 164.695 ;
        RECT 34.990 163.665 35.730 163.695 ;
        RECT 33.705 163.065 34.235 163.235 ;
        RECT 32.015 162.645 32.365 162.815 ;
        RECT 32.585 162.625 33.535 162.905 ;
        RECT 33.705 162.455 33.895 162.895 ;
        RECT 34.065 162.835 34.235 163.065 ;
        RECT 34.405 163.005 34.645 163.405 ;
        RECT 34.815 163.365 35.730 163.665 ;
        RECT 34.815 163.190 35.140 163.365 ;
        RECT 34.815 162.835 35.135 163.190 ;
        RECT 35.900 163.165 36.110 163.815 ;
        RECT 34.065 162.665 35.135 162.835 ;
        RECT 35.380 162.455 35.685 162.915 ;
        RECT 35.855 162.635 36.110 163.165 ;
        RECT 36.290 163.815 36.545 164.695 ;
        RECT 36.715 163.865 37.020 165.005 ;
        RECT 37.360 164.625 37.690 165.005 ;
        RECT 37.870 164.455 38.040 164.745 ;
        RECT 38.210 164.545 38.460 165.005 ;
        RECT 37.240 164.285 38.040 164.455 ;
        RECT 38.630 164.495 39.500 164.835 ;
        RECT 36.290 163.165 36.500 163.815 ;
        RECT 37.240 163.695 37.410 164.285 ;
        RECT 38.630 164.115 38.800 164.495 ;
        RECT 39.735 164.375 39.905 164.835 ;
        RECT 40.075 164.545 40.445 165.005 ;
        RECT 40.740 164.405 40.910 164.745 ;
        RECT 41.080 164.575 41.410 165.005 ;
        RECT 41.645 164.405 41.815 164.745 ;
        RECT 37.580 163.945 38.800 164.115 ;
        RECT 38.970 164.035 39.430 164.325 ;
        RECT 39.735 164.205 40.295 164.375 ;
        RECT 40.740 164.235 41.815 164.405 ;
        RECT 41.985 164.505 42.665 164.835 ;
        RECT 42.880 164.505 43.130 164.835 ;
        RECT 43.300 164.545 43.550 165.005 ;
        RECT 40.125 164.065 40.295 164.205 ;
        RECT 38.970 164.025 39.935 164.035 ;
        RECT 38.630 163.855 38.800 163.945 ;
        RECT 39.260 163.865 39.935 164.025 ;
        RECT 36.670 163.665 37.410 163.695 ;
        RECT 36.670 163.365 37.585 163.665 ;
        RECT 37.260 163.190 37.585 163.365 ;
        RECT 36.290 162.635 36.545 163.165 ;
        RECT 36.715 162.455 37.020 162.915 ;
        RECT 37.265 162.835 37.585 163.190 ;
        RECT 37.755 163.405 38.295 163.775 ;
        RECT 38.630 163.685 39.035 163.855 ;
        RECT 37.755 163.005 37.995 163.405 ;
        RECT 38.475 163.235 38.695 163.515 ;
        RECT 38.165 163.065 38.695 163.235 ;
        RECT 38.165 162.835 38.335 163.065 ;
        RECT 38.865 162.905 39.035 163.685 ;
        RECT 39.205 163.075 39.555 163.695 ;
        RECT 39.725 163.075 39.935 163.865 ;
        RECT 40.125 163.895 41.625 164.065 ;
        RECT 40.125 163.205 40.295 163.895 ;
        RECT 41.985 163.725 42.155 164.505 ;
        RECT 42.960 164.375 43.130 164.505 ;
        RECT 40.465 163.555 42.155 163.725 ;
        RECT 42.325 163.945 42.790 164.335 ;
        RECT 42.960 164.205 43.355 164.375 ;
        RECT 40.465 163.375 40.635 163.555 ;
        RECT 37.265 162.665 38.335 162.835 ;
        RECT 38.505 162.455 38.695 162.895 ;
        RECT 38.865 162.625 39.815 162.905 ;
        RECT 40.125 162.815 40.385 163.205 ;
        RECT 40.805 163.135 41.595 163.385 ;
        RECT 40.035 162.645 40.385 162.815 ;
        RECT 40.595 162.455 40.925 162.915 ;
        RECT 41.800 162.845 41.970 163.555 ;
        RECT 42.325 163.355 42.495 163.945 ;
        RECT 42.140 163.135 42.495 163.355 ;
        RECT 42.665 163.135 43.015 163.755 ;
        RECT 43.185 162.845 43.355 164.205 ;
        RECT 43.720 164.035 44.045 164.820 ;
        RECT 43.525 162.985 43.985 164.035 ;
        RECT 41.800 162.675 42.655 162.845 ;
        RECT 42.860 162.675 43.355 162.845 ;
        RECT 43.525 162.455 43.855 162.815 ;
        RECT 44.215 162.715 44.385 164.835 ;
        RECT 44.555 164.505 44.885 165.005 ;
        RECT 45.055 164.335 45.310 164.835 ;
        RECT 44.560 164.165 45.310 164.335 ;
        RECT 46.520 164.375 46.805 164.835 ;
        RECT 46.975 164.545 47.245 165.005 ;
        RECT 44.560 163.175 44.790 164.165 ;
        RECT 46.520 164.155 47.475 164.375 ;
        RECT 44.960 163.345 45.310 163.995 ;
        RECT 46.405 163.425 47.095 163.985 ;
        RECT 47.265 163.255 47.475 164.155 ;
        RECT 44.560 163.005 45.310 163.175 ;
        RECT 44.555 162.455 44.885 162.835 ;
        RECT 45.055 162.715 45.310 163.005 ;
        RECT 46.520 163.085 47.475 163.255 ;
        RECT 47.645 163.985 48.045 164.835 ;
        RECT 48.235 164.375 48.515 164.835 ;
        RECT 49.035 164.545 49.360 165.005 ;
        RECT 48.235 164.155 49.360 164.375 ;
        RECT 47.645 163.425 48.740 163.985 ;
        RECT 48.910 163.695 49.360 164.155 ;
        RECT 49.530 163.865 49.915 164.835 ;
        RECT 46.520 162.625 46.805 163.085 ;
        RECT 46.975 162.455 47.245 162.915 ;
        RECT 47.645 162.625 48.045 163.425 ;
        RECT 48.910 163.365 49.465 163.695 ;
        RECT 48.910 163.255 49.360 163.365 ;
        RECT 48.235 163.085 49.360 163.255 ;
        RECT 49.635 163.195 49.915 163.865 ;
        RECT 50.085 163.840 50.375 165.005 ;
        RECT 50.605 163.865 50.815 165.005 ;
        RECT 50.985 163.855 51.315 164.835 ;
        RECT 51.485 163.865 51.715 165.005 ;
        RECT 51.925 163.915 53.595 165.005 ;
        RECT 53.855 164.075 54.025 164.835 ;
        RECT 54.205 164.245 54.535 165.005 ;
        RECT 48.235 162.625 48.515 163.085 ;
        RECT 49.035 162.455 49.360 162.915 ;
        RECT 49.530 162.625 49.915 163.195 ;
        RECT 50.085 162.455 50.375 163.180 ;
        RECT 50.605 162.455 50.815 163.275 ;
        RECT 50.985 163.255 51.235 163.855 ;
        RECT 51.405 163.445 51.735 163.695 ;
        RECT 51.925 163.395 52.675 163.915 ;
        RECT 53.855 163.905 54.520 164.075 ;
        RECT 54.705 163.930 54.975 164.835 ;
        RECT 54.350 163.760 54.520 163.905 ;
        RECT 50.985 162.625 51.315 163.255 ;
        RECT 51.485 162.455 51.715 163.275 ;
        RECT 52.845 163.225 53.595 163.745 ;
        RECT 53.785 163.355 54.115 163.725 ;
        RECT 54.350 163.430 54.635 163.760 ;
        RECT 51.925 162.455 53.595 163.225 ;
        RECT 54.350 163.175 54.520 163.430 ;
        RECT 53.855 163.005 54.520 163.175 ;
        RECT 54.805 163.130 54.975 163.930 ;
        RECT 53.855 162.625 54.025 163.005 ;
        RECT 54.205 162.455 54.535 162.835 ;
        RECT 54.715 162.625 54.975 163.130 ;
        RECT 55.150 163.815 55.405 164.695 ;
        RECT 55.575 163.865 55.880 165.005 ;
        RECT 56.220 164.625 56.550 165.005 ;
        RECT 56.730 164.455 56.900 164.745 ;
        RECT 57.070 164.545 57.320 165.005 ;
        RECT 56.100 164.285 56.900 164.455 ;
        RECT 57.490 164.495 58.360 164.835 ;
        RECT 55.150 163.165 55.360 163.815 ;
        RECT 56.100 163.695 56.270 164.285 ;
        RECT 57.490 164.115 57.660 164.495 ;
        RECT 58.595 164.375 58.765 164.835 ;
        RECT 58.935 164.545 59.305 165.005 ;
        RECT 59.600 164.405 59.770 164.745 ;
        RECT 59.940 164.575 60.270 165.005 ;
        RECT 60.505 164.405 60.675 164.745 ;
        RECT 56.440 163.945 57.660 164.115 ;
        RECT 57.830 164.035 58.290 164.325 ;
        RECT 58.595 164.205 59.155 164.375 ;
        RECT 59.600 164.235 60.675 164.405 ;
        RECT 60.845 164.505 61.525 164.835 ;
        RECT 61.740 164.505 61.990 164.835 ;
        RECT 62.160 164.545 62.410 165.005 ;
        RECT 58.985 164.065 59.155 164.205 ;
        RECT 57.830 164.025 58.795 164.035 ;
        RECT 57.490 163.855 57.660 163.945 ;
        RECT 58.120 163.865 58.795 164.025 ;
        RECT 55.530 163.665 56.270 163.695 ;
        RECT 55.530 163.365 56.445 163.665 ;
        RECT 56.120 163.190 56.445 163.365 ;
        RECT 55.150 162.635 55.405 163.165 ;
        RECT 55.575 162.455 55.880 162.915 ;
        RECT 56.125 162.835 56.445 163.190 ;
        RECT 56.615 163.405 57.155 163.775 ;
        RECT 57.490 163.685 57.895 163.855 ;
        RECT 56.615 163.005 56.855 163.405 ;
        RECT 57.335 163.235 57.555 163.515 ;
        RECT 57.025 163.065 57.555 163.235 ;
        RECT 57.025 162.835 57.195 163.065 ;
        RECT 57.725 162.905 57.895 163.685 ;
        RECT 58.065 163.075 58.415 163.695 ;
        RECT 58.585 163.075 58.795 163.865 ;
        RECT 58.985 163.895 60.485 164.065 ;
        RECT 58.985 163.205 59.155 163.895 ;
        RECT 60.845 163.725 61.015 164.505 ;
        RECT 61.820 164.375 61.990 164.505 ;
        RECT 59.325 163.555 61.015 163.725 ;
        RECT 61.185 163.945 61.650 164.335 ;
        RECT 61.820 164.205 62.215 164.375 ;
        RECT 59.325 163.375 59.495 163.555 ;
        RECT 56.125 162.665 57.195 162.835 ;
        RECT 57.365 162.455 57.555 162.895 ;
        RECT 57.725 162.625 58.675 162.905 ;
        RECT 58.985 162.815 59.245 163.205 ;
        RECT 59.665 163.135 60.455 163.385 ;
        RECT 58.895 162.645 59.245 162.815 ;
        RECT 59.455 162.455 59.785 162.915 ;
        RECT 60.660 162.845 60.830 163.555 ;
        RECT 61.185 163.355 61.355 163.945 ;
        RECT 61.000 163.135 61.355 163.355 ;
        RECT 61.525 163.135 61.875 163.755 ;
        RECT 62.045 162.845 62.215 164.205 ;
        RECT 62.580 164.035 62.905 164.820 ;
        RECT 62.385 162.985 62.845 164.035 ;
        RECT 60.660 162.675 61.515 162.845 ;
        RECT 61.720 162.675 62.215 162.845 ;
        RECT 62.385 162.455 62.715 162.815 ;
        RECT 63.075 162.715 63.245 164.835 ;
        RECT 63.415 164.505 63.745 165.005 ;
        RECT 63.915 164.335 64.170 164.835 ;
        RECT 63.420 164.165 64.170 164.335 ;
        RECT 63.420 163.175 63.650 164.165 ;
        RECT 63.820 163.345 64.170 163.995 ;
        RECT 64.495 163.855 64.825 165.005 ;
        RECT 64.995 163.985 65.165 164.835 ;
        RECT 65.335 164.205 65.665 165.005 ;
        RECT 65.835 163.985 66.005 164.835 ;
        RECT 66.185 164.205 66.425 165.005 ;
        RECT 66.595 164.025 66.925 164.835 ;
        RECT 67.160 164.135 67.445 165.005 ;
        RECT 67.615 164.375 67.875 164.835 ;
        RECT 68.050 164.545 68.305 165.005 ;
        RECT 68.475 164.375 68.735 164.835 ;
        RECT 67.615 164.205 68.735 164.375 ;
        RECT 68.905 164.205 69.215 165.005 ;
        RECT 64.995 163.815 66.005 163.985 ;
        RECT 66.210 163.855 66.925 164.025 ;
        RECT 67.615 163.955 67.875 164.205 ;
        RECT 69.385 164.035 69.695 164.835 ;
        RECT 70.330 164.570 75.675 165.005 ;
        RECT 64.995 163.305 65.490 163.815 ;
        RECT 66.210 163.615 66.380 163.855 ;
        RECT 67.120 163.785 67.875 163.955 ;
        RECT 68.665 163.865 69.695 164.035 ;
        RECT 65.880 163.445 66.380 163.615 ;
        RECT 66.550 163.445 66.930 163.685 ;
        RECT 64.995 163.275 65.495 163.305 ;
        RECT 66.210 163.275 66.380 163.445 ;
        RECT 67.120 163.275 67.525 163.785 ;
        RECT 68.665 163.615 68.835 163.865 ;
        RECT 67.695 163.445 68.835 163.615 ;
        RECT 63.420 163.005 64.170 163.175 ;
        RECT 63.415 162.455 63.745 162.835 ;
        RECT 63.915 162.715 64.170 163.005 ;
        RECT 64.495 162.455 64.825 163.255 ;
        RECT 64.995 163.105 66.005 163.275 ;
        RECT 66.210 163.105 66.845 163.275 ;
        RECT 67.120 163.105 68.770 163.275 ;
        RECT 69.005 163.125 69.355 163.695 ;
        RECT 64.995 162.625 65.165 163.105 ;
        RECT 65.335 162.455 65.665 162.935 ;
        RECT 65.835 162.625 66.005 163.105 ;
        RECT 66.255 162.455 66.495 162.935 ;
        RECT 66.675 162.625 66.845 163.105 ;
        RECT 67.165 162.455 67.445 162.935 ;
        RECT 67.615 162.715 67.875 163.105 ;
        RECT 68.050 162.455 68.305 162.935 ;
        RECT 68.475 162.715 68.770 163.105 ;
        RECT 69.525 162.955 69.695 163.865 ;
        RECT 71.920 163.320 72.270 164.570 ;
        RECT 75.845 163.840 76.135 165.005 ;
        RECT 76.305 163.915 77.975 165.005 ;
        RECT 78.145 164.245 78.660 164.655 ;
        RECT 78.895 164.245 79.065 165.005 ;
        RECT 79.235 164.665 81.265 164.835 ;
        RECT 73.750 163.000 74.090 163.830 ;
        RECT 76.305 163.395 77.055 163.915 ;
        RECT 77.225 163.225 77.975 163.745 ;
        RECT 78.145 163.435 78.485 164.245 ;
        RECT 79.235 164.000 79.405 164.665 ;
        RECT 79.800 164.325 80.925 164.495 ;
        RECT 78.655 163.810 79.405 164.000 ;
        RECT 79.575 163.985 80.585 164.155 ;
        RECT 78.145 163.265 79.375 163.435 ;
        RECT 68.950 162.455 69.225 162.935 ;
        RECT 69.395 162.625 69.695 162.955 ;
        RECT 70.330 162.455 75.675 163.000 ;
        RECT 75.845 162.455 76.135 163.180 ;
        RECT 76.305 162.455 77.975 163.225 ;
        RECT 78.420 162.660 78.665 163.265 ;
        RECT 78.885 162.455 79.395 162.990 ;
        RECT 79.575 162.625 79.765 163.985 ;
        RECT 79.935 162.965 80.210 163.785 ;
        RECT 80.415 163.185 80.585 163.985 ;
        RECT 80.755 163.195 80.925 164.325 ;
        RECT 81.095 163.695 81.265 164.665 ;
        RECT 81.435 163.865 81.605 165.005 ;
        RECT 81.775 163.865 82.110 164.835 ;
        RECT 82.375 164.075 82.545 164.835 ;
        RECT 82.725 164.245 83.055 165.005 ;
        RECT 82.375 163.905 83.040 164.075 ;
        RECT 83.225 163.930 83.495 164.835 ;
        RECT 81.095 163.365 81.290 163.695 ;
        RECT 81.515 163.365 81.770 163.695 ;
        RECT 81.515 163.195 81.685 163.365 ;
        RECT 81.940 163.195 82.110 163.865 ;
        RECT 82.870 163.760 83.040 163.905 ;
        RECT 82.305 163.355 82.635 163.725 ;
        RECT 82.870 163.430 83.155 163.760 ;
        RECT 80.755 163.025 81.685 163.195 ;
        RECT 80.755 162.990 80.930 163.025 ;
        RECT 79.935 162.795 80.215 162.965 ;
        RECT 79.935 162.625 80.210 162.795 ;
        RECT 80.400 162.625 80.930 162.990 ;
        RECT 81.355 162.455 81.685 162.855 ;
        RECT 81.855 162.625 82.110 163.195 ;
        RECT 82.870 163.175 83.040 163.430 ;
        RECT 82.375 163.005 83.040 163.175 ;
        RECT 83.325 163.130 83.495 163.930 ;
        RECT 83.665 163.915 85.335 165.005 ;
        RECT 85.595 164.075 85.765 164.835 ;
        RECT 85.945 164.245 86.275 165.005 ;
        RECT 83.665 163.395 84.415 163.915 ;
        RECT 85.595 163.905 86.260 164.075 ;
        RECT 86.445 163.930 86.715 164.835 ;
        RECT 86.890 164.570 92.235 165.005 ;
        RECT 86.090 163.760 86.260 163.905 ;
        RECT 84.585 163.225 85.335 163.745 ;
        RECT 85.525 163.355 85.855 163.725 ;
        RECT 86.090 163.430 86.375 163.760 ;
        RECT 82.375 162.625 82.545 163.005 ;
        RECT 82.725 162.455 83.055 162.835 ;
        RECT 83.235 162.625 83.495 163.130 ;
        RECT 83.665 162.455 85.335 163.225 ;
        RECT 86.090 163.175 86.260 163.430 ;
        RECT 85.595 163.005 86.260 163.175 ;
        RECT 86.545 163.130 86.715 163.930 ;
        RECT 88.480 163.320 88.830 164.570 ;
        RECT 92.495 164.260 92.765 165.005 ;
        RECT 93.395 165.000 99.670 165.005 ;
        RECT 92.935 164.090 93.225 164.830 ;
        RECT 93.395 164.275 93.650 165.000 ;
        RECT 93.835 164.105 94.095 164.830 ;
        RECT 94.265 164.275 94.510 165.000 ;
        RECT 94.695 164.105 94.955 164.830 ;
        RECT 95.125 164.275 95.370 165.000 ;
        RECT 95.555 164.105 95.815 164.830 ;
        RECT 95.985 164.275 96.230 165.000 ;
        RECT 96.400 164.105 96.660 164.830 ;
        RECT 96.830 164.275 97.090 165.000 ;
        RECT 97.260 164.105 97.520 164.830 ;
        RECT 97.690 164.275 97.950 165.000 ;
        RECT 98.120 164.105 98.380 164.830 ;
        RECT 98.550 164.275 98.810 165.000 ;
        RECT 98.980 164.105 99.240 164.830 ;
        RECT 99.410 164.205 99.670 165.000 ;
        RECT 93.835 164.090 99.240 164.105 ;
        RECT 92.495 163.865 99.240 164.090 ;
        RECT 85.595 162.625 85.765 163.005 ;
        RECT 85.945 162.455 86.275 162.835 ;
        RECT 86.455 162.625 86.715 163.130 ;
        RECT 90.310 163.000 90.650 163.830 ;
        RECT 92.495 163.275 93.660 163.865 ;
        RECT 99.840 163.695 100.090 164.830 ;
        RECT 100.270 164.195 100.530 165.005 ;
        RECT 100.705 163.695 100.950 164.835 ;
        RECT 101.130 164.195 101.425 165.005 ;
        RECT 101.605 163.840 101.895 165.005 ;
        RECT 102.065 164.245 102.580 164.655 ;
        RECT 102.815 164.245 102.985 165.005 ;
        RECT 103.155 164.665 105.185 164.835 ;
        RECT 93.830 163.445 100.950 163.695 ;
        RECT 92.495 163.105 99.240 163.275 ;
        RECT 86.890 162.455 92.235 163.000 ;
        RECT 92.495 162.455 92.795 162.935 ;
        RECT 92.965 162.650 93.225 163.105 ;
        RECT 93.395 162.455 93.655 162.935 ;
        RECT 93.835 162.650 94.095 163.105 ;
        RECT 94.265 162.455 94.515 162.935 ;
        RECT 94.695 162.650 94.955 163.105 ;
        RECT 95.125 162.455 95.375 162.935 ;
        RECT 95.555 162.650 95.815 163.105 ;
        RECT 95.985 162.455 96.230 162.935 ;
        RECT 96.400 162.650 96.675 163.105 ;
        RECT 96.845 162.455 97.090 162.935 ;
        RECT 97.260 162.650 97.520 163.105 ;
        RECT 97.690 162.455 97.950 162.935 ;
        RECT 98.120 162.650 98.380 163.105 ;
        RECT 98.550 162.455 98.810 162.935 ;
        RECT 98.980 162.650 99.240 163.105 ;
        RECT 99.410 162.455 99.670 163.015 ;
        RECT 99.840 162.635 100.090 163.445 ;
        RECT 100.270 162.455 100.530 162.980 ;
        RECT 100.700 162.635 100.950 163.445 ;
        RECT 101.120 163.135 101.435 163.695 ;
        RECT 102.065 163.435 102.405 164.245 ;
        RECT 103.155 164.000 103.325 164.665 ;
        RECT 103.720 164.325 104.845 164.495 ;
        RECT 102.575 163.810 103.325 164.000 ;
        RECT 103.495 163.985 104.505 164.155 ;
        RECT 102.065 163.265 103.295 163.435 ;
        RECT 101.130 162.455 101.435 162.965 ;
        RECT 101.605 162.455 101.895 163.180 ;
        RECT 102.340 162.660 102.585 163.265 ;
        RECT 102.805 162.455 103.315 162.990 ;
        RECT 103.495 162.625 103.685 163.985 ;
        RECT 103.855 163.305 104.130 163.785 ;
        RECT 103.855 163.135 104.135 163.305 ;
        RECT 104.335 163.185 104.505 163.985 ;
        RECT 104.675 163.195 104.845 164.325 ;
        RECT 105.015 163.695 105.185 164.665 ;
        RECT 105.355 163.865 105.525 165.005 ;
        RECT 105.695 163.865 106.030 164.835 ;
        RECT 105.015 163.365 105.210 163.695 ;
        RECT 105.435 163.365 105.690 163.695 ;
        RECT 105.435 163.195 105.605 163.365 ;
        RECT 105.860 163.195 106.030 163.865 ;
        RECT 103.855 162.625 104.130 163.135 ;
        RECT 104.675 163.025 105.605 163.195 ;
        RECT 104.675 162.990 104.850 163.025 ;
        RECT 104.320 162.625 104.850 162.990 ;
        RECT 105.275 162.455 105.605 162.855 ;
        RECT 105.775 162.625 106.030 163.195 ;
        RECT 106.670 163.865 107.005 164.835 ;
        RECT 107.175 163.865 107.345 165.005 ;
        RECT 107.515 164.665 109.545 164.835 ;
        RECT 106.670 163.195 106.840 163.865 ;
        RECT 107.515 163.695 107.685 164.665 ;
        RECT 107.010 163.365 107.265 163.695 ;
        RECT 107.490 163.365 107.685 163.695 ;
        RECT 107.855 164.325 108.980 164.495 ;
        RECT 107.095 163.195 107.265 163.365 ;
        RECT 107.855 163.195 108.025 164.325 ;
        RECT 106.670 162.625 106.925 163.195 ;
        RECT 107.095 163.025 108.025 163.195 ;
        RECT 108.195 163.985 109.205 164.155 ;
        RECT 108.195 163.185 108.365 163.985 ;
        RECT 107.850 162.990 108.025 163.025 ;
        RECT 107.095 162.455 107.425 162.855 ;
        RECT 107.850 162.625 108.380 162.990 ;
        RECT 108.570 162.965 108.845 163.785 ;
        RECT 108.565 162.795 108.845 162.965 ;
        RECT 108.570 162.625 108.845 162.795 ;
        RECT 109.015 162.625 109.205 163.985 ;
        RECT 109.375 164.000 109.545 164.665 ;
        RECT 109.715 164.245 109.885 165.005 ;
        RECT 110.120 164.245 110.635 164.655 ;
        RECT 109.375 163.810 110.125 164.000 ;
        RECT 110.295 163.435 110.635 164.245 ;
        RECT 110.955 163.855 111.285 165.005 ;
        RECT 111.455 163.985 111.625 164.835 ;
        RECT 111.795 164.205 112.125 165.005 ;
        RECT 112.295 163.985 112.465 164.835 ;
        RECT 112.645 164.205 112.885 165.005 ;
        RECT 113.055 164.025 113.385 164.835 ;
        RECT 109.405 163.265 110.635 163.435 ;
        RECT 111.455 163.815 112.465 163.985 ;
        RECT 112.670 163.855 113.385 164.025 ;
        RECT 111.455 163.305 111.950 163.815 ;
        RECT 112.670 163.615 112.840 163.855 ;
        RECT 113.570 163.815 113.825 164.695 ;
        RECT 113.995 163.865 114.300 165.005 ;
        RECT 114.640 164.625 114.970 165.005 ;
        RECT 115.150 164.455 115.320 164.745 ;
        RECT 115.490 164.545 115.740 165.005 ;
        RECT 114.520 164.285 115.320 164.455 ;
        RECT 115.910 164.495 116.780 164.835 ;
        RECT 112.340 163.445 112.840 163.615 ;
        RECT 113.010 163.445 113.390 163.685 ;
        RECT 111.455 163.275 111.955 163.305 ;
        RECT 112.670 163.275 112.840 163.445 ;
        RECT 109.385 162.455 109.895 162.990 ;
        RECT 110.115 162.660 110.360 163.265 ;
        RECT 110.955 162.455 111.285 163.255 ;
        RECT 111.455 163.105 112.465 163.275 ;
        RECT 112.670 163.105 113.305 163.275 ;
        RECT 111.455 162.625 111.625 163.105 ;
        RECT 111.795 162.455 112.125 162.935 ;
        RECT 112.295 162.625 112.465 163.105 ;
        RECT 112.715 162.455 112.955 162.935 ;
        RECT 113.135 162.625 113.305 163.105 ;
        RECT 113.570 163.165 113.780 163.815 ;
        RECT 114.520 163.695 114.690 164.285 ;
        RECT 115.910 164.115 116.080 164.495 ;
        RECT 117.015 164.375 117.185 164.835 ;
        RECT 117.355 164.545 117.725 165.005 ;
        RECT 118.020 164.405 118.190 164.745 ;
        RECT 118.360 164.575 118.690 165.005 ;
        RECT 118.925 164.405 119.095 164.745 ;
        RECT 114.860 163.945 116.080 164.115 ;
        RECT 116.250 164.035 116.710 164.325 ;
        RECT 117.015 164.205 117.575 164.375 ;
        RECT 118.020 164.235 119.095 164.405 ;
        RECT 119.265 164.505 119.945 164.835 ;
        RECT 120.160 164.505 120.410 164.835 ;
        RECT 120.580 164.545 120.830 165.005 ;
        RECT 117.405 164.065 117.575 164.205 ;
        RECT 116.250 164.025 117.215 164.035 ;
        RECT 115.910 163.855 116.080 163.945 ;
        RECT 116.540 163.865 117.215 164.025 ;
        RECT 113.950 163.665 114.690 163.695 ;
        RECT 113.950 163.365 114.865 163.665 ;
        RECT 114.540 163.190 114.865 163.365 ;
        RECT 113.570 162.635 113.825 163.165 ;
        RECT 113.995 162.455 114.300 162.915 ;
        RECT 114.545 162.835 114.865 163.190 ;
        RECT 115.035 163.405 115.575 163.775 ;
        RECT 115.910 163.685 116.315 163.855 ;
        RECT 115.035 163.005 115.275 163.405 ;
        RECT 115.755 163.235 115.975 163.515 ;
        RECT 115.445 163.065 115.975 163.235 ;
        RECT 115.445 162.835 115.615 163.065 ;
        RECT 116.145 162.905 116.315 163.685 ;
        RECT 116.485 163.075 116.835 163.695 ;
        RECT 117.005 163.075 117.215 163.865 ;
        RECT 117.405 163.895 118.905 164.065 ;
        RECT 117.405 163.205 117.575 163.895 ;
        RECT 119.265 163.725 119.435 164.505 ;
        RECT 120.240 164.375 120.410 164.505 ;
        RECT 117.745 163.555 119.435 163.725 ;
        RECT 119.605 163.945 120.070 164.335 ;
        RECT 120.240 164.205 120.635 164.375 ;
        RECT 117.745 163.375 117.915 163.555 ;
        RECT 114.545 162.665 115.615 162.835 ;
        RECT 115.785 162.455 115.975 162.895 ;
        RECT 116.145 162.625 117.095 162.905 ;
        RECT 117.405 162.815 117.665 163.205 ;
        RECT 118.085 163.135 118.875 163.385 ;
        RECT 117.315 162.645 117.665 162.815 ;
        RECT 117.875 162.455 118.205 162.915 ;
        RECT 119.080 162.845 119.250 163.555 ;
        RECT 119.605 163.355 119.775 163.945 ;
        RECT 119.420 163.135 119.775 163.355 ;
        RECT 119.945 163.135 120.295 163.755 ;
        RECT 120.465 162.845 120.635 164.205 ;
        RECT 121.000 164.035 121.325 164.820 ;
        RECT 120.805 162.985 121.265 164.035 ;
        RECT 119.080 162.675 119.935 162.845 ;
        RECT 120.140 162.675 120.635 162.845 ;
        RECT 120.805 162.455 121.135 162.815 ;
        RECT 121.495 162.715 121.665 164.835 ;
        RECT 121.835 164.505 122.165 165.005 ;
        RECT 122.335 164.335 122.590 164.835 ;
        RECT 121.840 164.165 122.590 164.335 ;
        RECT 121.840 163.175 122.070 164.165 ;
        RECT 122.240 163.345 122.590 163.995 ;
        RECT 122.765 163.930 123.035 164.835 ;
        RECT 123.205 164.245 123.535 165.005 ;
        RECT 123.715 164.075 123.885 164.835 ;
        RECT 121.840 163.005 122.590 163.175 ;
        RECT 121.835 162.455 122.165 162.835 ;
        RECT 122.335 162.715 122.590 163.005 ;
        RECT 122.765 163.130 122.935 163.930 ;
        RECT 123.220 163.905 123.885 164.075 ;
        RECT 124.605 163.915 126.275 165.005 ;
        RECT 126.445 163.915 127.655 165.005 ;
        RECT 123.220 163.760 123.390 163.905 ;
        RECT 123.105 163.430 123.390 163.760 ;
        RECT 123.220 163.175 123.390 163.430 ;
        RECT 123.625 163.355 123.955 163.725 ;
        RECT 124.605 163.395 125.355 163.915 ;
        RECT 125.525 163.225 126.275 163.745 ;
        RECT 126.445 163.375 126.965 163.915 ;
        RECT 122.765 162.625 123.025 163.130 ;
        RECT 123.220 163.005 123.885 163.175 ;
        RECT 123.205 162.455 123.535 162.835 ;
        RECT 123.715 162.625 123.885 163.005 ;
        RECT 124.605 162.455 126.275 163.225 ;
        RECT 127.135 163.205 127.655 163.745 ;
        RECT 126.445 162.455 127.655 163.205 ;
        RECT 14.580 162.285 127.740 162.455 ;
        RECT 14.665 161.535 15.875 162.285 ;
        RECT 14.665 160.995 15.185 161.535 ;
        RECT 16.045 161.515 17.715 162.285 ;
        RECT 15.355 160.825 15.875 161.365 ;
        RECT 14.665 159.735 15.875 160.825 ;
        RECT 16.045 160.825 16.795 161.345 ;
        RECT 16.965 160.995 17.715 161.515 ;
        RECT 18.260 161.575 18.515 162.105 ;
        RECT 18.695 161.825 18.980 162.285 ;
        RECT 16.045 159.735 17.715 160.825 ;
        RECT 18.260 160.715 18.440 161.575 ;
        RECT 19.160 161.375 19.410 162.025 ;
        RECT 18.610 161.045 19.410 161.375 ;
        RECT 18.260 160.245 18.515 160.715 ;
        RECT 18.175 160.075 18.515 160.245 ;
        RECT 18.260 160.045 18.515 160.075 ;
        RECT 18.695 159.735 18.980 160.535 ;
        RECT 19.160 160.455 19.410 161.045 ;
        RECT 19.610 161.690 19.930 162.020 ;
        RECT 20.110 161.805 20.770 162.285 ;
        RECT 20.970 161.895 21.820 162.065 ;
        RECT 19.610 160.795 19.800 161.690 ;
        RECT 20.120 161.365 20.780 161.635 ;
        RECT 20.450 161.305 20.780 161.365 ;
        RECT 19.970 161.135 20.300 161.195 ;
        RECT 20.970 161.135 21.140 161.895 ;
        RECT 22.380 161.825 22.700 162.285 ;
        RECT 22.900 161.645 23.150 162.075 ;
        RECT 23.440 161.845 23.850 162.285 ;
        RECT 24.020 161.905 25.035 162.105 ;
        RECT 21.310 161.475 22.560 161.645 ;
        RECT 21.310 161.355 21.640 161.475 ;
        RECT 19.970 160.965 21.870 161.135 ;
        RECT 19.610 160.625 21.530 160.795 ;
        RECT 19.610 160.605 19.930 160.625 ;
        RECT 19.160 159.945 19.490 160.455 ;
        RECT 19.760 159.995 19.930 160.605 ;
        RECT 21.700 160.455 21.870 160.965 ;
        RECT 22.040 160.895 22.220 161.305 ;
        RECT 22.390 160.715 22.560 161.475 ;
        RECT 20.100 159.735 20.430 160.425 ;
        RECT 20.660 160.285 21.870 160.455 ;
        RECT 22.040 160.405 22.560 160.715 ;
        RECT 22.730 161.305 23.150 161.645 ;
        RECT 23.440 161.305 23.850 161.635 ;
        RECT 22.730 160.535 22.920 161.305 ;
        RECT 24.020 161.175 24.190 161.905 ;
        RECT 25.335 161.735 25.505 162.065 ;
        RECT 25.675 161.905 26.005 162.285 ;
        RECT 24.360 161.355 24.710 161.725 ;
        RECT 24.020 161.135 24.440 161.175 ;
        RECT 23.090 160.965 24.440 161.135 ;
        RECT 23.090 160.805 23.340 160.965 ;
        RECT 23.850 160.535 24.100 160.795 ;
        RECT 22.730 160.285 24.100 160.535 ;
        RECT 20.660 159.995 20.900 160.285 ;
        RECT 21.700 160.205 21.870 160.285 ;
        RECT 21.100 159.735 21.520 160.115 ;
        RECT 21.700 159.955 22.330 160.205 ;
        RECT 22.800 159.735 23.130 160.115 ;
        RECT 23.300 159.995 23.470 160.285 ;
        RECT 24.270 160.120 24.440 160.965 ;
        RECT 24.890 160.795 25.110 161.665 ;
        RECT 25.335 161.545 26.030 161.735 ;
        RECT 24.610 160.415 25.110 160.795 ;
        RECT 25.280 160.745 25.690 161.365 ;
        RECT 25.860 160.575 26.030 161.545 ;
        RECT 25.335 160.405 26.030 160.575 ;
        RECT 23.650 159.735 24.030 160.115 ;
        RECT 24.270 159.950 25.100 160.120 ;
        RECT 25.335 159.905 25.505 160.405 ;
        RECT 25.675 159.735 26.005 160.235 ;
        RECT 26.220 159.905 26.445 162.025 ;
        RECT 26.615 161.905 26.945 162.285 ;
        RECT 27.115 161.735 27.285 162.025 ;
        RECT 26.620 161.565 27.285 161.735 ;
        RECT 26.620 160.575 26.850 161.565 ;
        RECT 27.550 161.545 27.805 162.115 ;
        RECT 27.975 161.885 28.305 162.285 ;
        RECT 28.730 161.750 29.260 162.115 ;
        RECT 28.730 161.715 28.905 161.750 ;
        RECT 27.975 161.545 28.905 161.715 ;
        RECT 29.450 161.605 29.725 162.115 ;
        RECT 27.020 160.745 27.370 161.395 ;
        RECT 27.550 160.875 27.720 161.545 ;
        RECT 27.975 161.375 28.145 161.545 ;
        RECT 27.890 161.045 28.145 161.375 ;
        RECT 28.370 161.045 28.565 161.375 ;
        RECT 26.620 160.405 27.285 160.575 ;
        RECT 26.615 159.735 26.945 160.235 ;
        RECT 27.115 159.905 27.285 160.405 ;
        RECT 27.550 159.905 27.885 160.875 ;
        RECT 28.055 159.735 28.225 160.875 ;
        RECT 28.395 160.075 28.565 161.045 ;
        RECT 28.735 160.415 28.905 161.545 ;
        RECT 29.075 160.755 29.245 161.555 ;
        RECT 29.445 161.435 29.725 161.605 ;
        RECT 29.450 160.955 29.725 161.435 ;
        RECT 29.895 160.755 30.085 162.115 ;
        RECT 30.265 161.750 30.775 162.285 ;
        RECT 30.995 161.475 31.240 162.080 ;
        RECT 31.685 161.535 32.895 162.285 ;
        RECT 30.285 161.305 31.515 161.475 ;
        RECT 29.075 160.585 30.085 160.755 ;
        RECT 30.255 160.740 31.005 160.930 ;
        RECT 28.735 160.245 29.860 160.415 ;
        RECT 30.255 160.075 30.425 160.740 ;
        RECT 31.175 160.495 31.515 161.305 ;
        RECT 28.395 159.905 30.425 160.075 ;
        RECT 30.595 159.735 30.765 160.495 ;
        RECT 31.000 160.085 31.515 160.495 ;
        RECT 31.685 160.825 32.205 161.365 ;
        RECT 32.375 160.995 32.895 161.535 ;
        RECT 33.070 161.545 33.325 162.115 ;
        RECT 33.495 161.885 33.825 162.285 ;
        RECT 34.250 161.750 34.780 162.115 ;
        RECT 34.250 161.715 34.425 161.750 ;
        RECT 33.495 161.545 34.425 161.715 ;
        RECT 34.970 161.605 35.245 162.115 ;
        RECT 33.070 160.875 33.240 161.545 ;
        RECT 33.495 161.375 33.665 161.545 ;
        RECT 33.410 161.045 33.665 161.375 ;
        RECT 33.890 161.045 34.085 161.375 ;
        RECT 31.685 159.735 32.895 160.825 ;
        RECT 33.070 159.905 33.405 160.875 ;
        RECT 33.575 159.735 33.745 160.875 ;
        RECT 33.915 160.075 34.085 161.045 ;
        RECT 34.255 160.415 34.425 161.545 ;
        RECT 34.595 160.755 34.765 161.555 ;
        RECT 34.965 161.435 35.245 161.605 ;
        RECT 34.970 160.955 35.245 161.435 ;
        RECT 35.415 160.755 35.605 162.115 ;
        RECT 35.785 161.750 36.295 162.285 ;
        RECT 36.515 161.475 36.760 162.080 ;
        RECT 37.205 161.560 37.495 162.285 ;
        RECT 38.125 161.515 39.795 162.285 ;
        RECT 35.805 161.305 37.035 161.475 ;
        RECT 34.595 160.585 35.605 160.755 ;
        RECT 35.775 160.740 36.525 160.930 ;
        RECT 34.255 160.245 35.380 160.415 ;
        RECT 35.775 160.075 35.945 160.740 ;
        RECT 36.695 160.495 37.035 161.305 ;
        RECT 33.915 159.905 35.945 160.075 ;
        RECT 36.115 159.735 36.285 160.495 ;
        RECT 36.520 160.085 37.035 160.495 ;
        RECT 37.205 159.735 37.495 160.900 ;
        RECT 38.125 160.825 38.875 161.345 ;
        RECT 39.045 160.995 39.795 161.515 ;
        RECT 40.080 161.655 40.365 162.115 ;
        RECT 40.535 161.825 40.805 162.285 ;
        RECT 40.080 161.485 41.035 161.655 ;
        RECT 38.125 159.735 39.795 160.825 ;
        RECT 39.965 160.755 40.655 161.315 ;
        RECT 40.825 160.585 41.035 161.485 ;
        RECT 40.080 160.365 41.035 160.585 ;
        RECT 41.205 161.315 41.605 162.115 ;
        RECT 41.795 161.655 42.075 162.115 ;
        RECT 42.595 161.825 42.920 162.285 ;
        RECT 41.795 161.485 42.920 161.655 ;
        RECT 43.090 161.545 43.475 162.115 ;
        RECT 42.470 161.375 42.920 161.485 ;
        RECT 41.205 160.755 42.300 161.315 ;
        RECT 42.470 161.045 43.025 161.375 ;
        RECT 40.080 159.905 40.365 160.365 ;
        RECT 40.535 159.735 40.805 160.195 ;
        RECT 41.205 159.905 41.605 160.755 ;
        RECT 42.470 160.585 42.920 161.045 ;
        RECT 43.195 160.875 43.475 161.545 ;
        RECT 41.795 160.365 42.920 160.585 ;
        RECT 41.795 159.905 42.075 160.365 ;
        RECT 42.595 159.735 42.920 160.195 ;
        RECT 43.090 159.905 43.475 160.875 ;
        RECT 43.650 161.545 43.905 162.115 ;
        RECT 44.075 161.885 44.405 162.285 ;
        RECT 44.830 161.750 45.360 162.115 ;
        RECT 45.550 161.945 45.825 162.115 ;
        RECT 45.545 161.775 45.825 161.945 ;
        RECT 44.830 161.715 45.005 161.750 ;
        RECT 44.075 161.545 45.005 161.715 ;
        RECT 43.650 160.875 43.820 161.545 ;
        RECT 44.075 161.375 44.245 161.545 ;
        RECT 43.990 161.045 44.245 161.375 ;
        RECT 44.470 161.045 44.665 161.375 ;
        RECT 43.650 159.905 43.985 160.875 ;
        RECT 44.155 159.735 44.325 160.875 ;
        RECT 44.495 160.075 44.665 161.045 ;
        RECT 44.835 160.415 45.005 161.545 ;
        RECT 45.175 160.755 45.345 161.555 ;
        RECT 45.550 160.955 45.825 161.775 ;
        RECT 45.995 160.755 46.185 162.115 ;
        RECT 46.365 161.750 46.875 162.285 ;
        RECT 47.095 161.475 47.340 162.080 ;
        RECT 47.785 161.610 48.045 162.115 ;
        RECT 48.225 161.905 48.555 162.285 ;
        RECT 48.735 161.735 48.905 162.115 ;
        RECT 46.385 161.305 47.615 161.475 ;
        RECT 45.175 160.585 46.185 160.755 ;
        RECT 46.355 160.740 47.105 160.930 ;
        RECT 44.835 160.245 45.960 160.415 ;
        RECT 46.355 160.075 46.525 160.740 ;
        RECT 47.275 160.495 47.615 161.305 ;
        RECT 44.495 159.905 46.525 160.075 ;
        RECT 46.695 159.735 46.865 160.495 ;
        RECT 47.100 160.085 47.615 160.495 ;
        RECT 47.785 160.810 47.955 161.610 ;
        RECT 48.240 161.565 48.905 161.735 ;
        RECT 48.240 161.310 48.410 161.565 ;
        RECT 49.170 161.545 49.425 162.115 ;
        RECT 49.595 161.885 49.925 162.285 ;
        RECT 50.350 161.750 50.880 162.115 ;
        RECT 50.350 161.715 50.525 161.750 ;
        RECT 49.595 161.545 50.525 161.715 ;
        RECT 48.125 160.980 48.410 161.310 ;
        RECT 48.645 161.015 48.975 161.385 ;
        RECT 48.240 160.835 48.410 160.980 ;
        RECT 49.170 160.875 49.340 161.545 ;
        RECT 49.595 161.375 49.765 161.545 ;
        RECT 49.510 161.045 49.765 161.375 ;
        RECT 49.990 161.045 50.185 161.375 ;
        RECT 47.785 159.905 48.055 160.810 ;
        RECT 48.240 160.665 48.905 160.835 ;
        RECT 48.225 159.735 48.555 160.495 ;
        RECT 48.735 159.905 48.905 160.665 ;
        RECT 49.170 159.905 49.505 160.875 ;
        RECT 49.675 159.735 49.845 160.875 ;
        RECT 50.015 160.075 50.185 161.045 ;
        RECT 50.355 160.415 50.525 161.545 ;
        RECT 50.695 160.755 50.865 161.555 ;
        RECT 51.070 161.265 51.345 162.115 ;
        RECT 51.065 161.095 51.345 161.265 ;
        RECT 51.070 160.955 51.345 161.095 ;
        RECT 51.515 160.755 51.705 162.115 ;
        RECT 51.885 161.750 52.395 162.285 ;
        RECT 52.615 161.475 52.860 162.080 ;
        RECT 53.580 161.475 53.825 162.080 ;
        RECT 54.045 161.750 54.555 162.285 ;
        RECT 51.905 161.305 53.135 161.475 ;
        RECT 50.695 160.585 51.705 160.755 ;
        RECT 51.875 160.740 52.625 160.930 ;
        RECT 50.355 160.245 51.480 160.415 ;
        RECT 51.875 160.075 52.045 160.740 ;
        RECT 52.795 160.495 53.135 161.305 ;
        RECT 50.015 159.905 52.045 160.075 ;
        RECT 52.215 159.735 52.385 160.495 ;
        RECT 52.620 160.085 53.135 160.495 ;
        RECT 53.305 161.305 54.535 161.475 ;
        RECT 53.305 160.495 53.645 161.305 ;
        RECT 53.815 160.740 54.565 160.930 ;
        RECT 53.305 160.085 53.820 160.495 ;
        RECT 54.055 159.735 54.225 160.495 ;
        RECT 54.395 160.075 54.565 160.740 ;
        RECT 54.735 160.755 54.925 162.115 ;
        RECT 55.095 161.945 55.370 162.115 ;
        RECT 55.095 161.775 55.375 161.945 ;
        RECT 55.095 160.955 55.370 161.775 ;
        RECT 55.560 161.750 56.090 162.115 ;
        RECT 56.515 161.885 56.845 162.285 ;
        RECT 55.915 161.715 56.090 161.750 ;
        RECT 55.575 160.755 55.745 161.555 ;
        RECT 54.735 160.585 55.745 160.755 ;
        RECT 55.915 161.545 56.845 161.715 ;
        RECT 57.015 161.545 57.270 162.115 ;
        RECT 55.915 160.415 56.085 161.545 ;
        RECT 56.675 161.375 56.845 161.545 ;
        RECT 54.960 160.245 56.085 160.415 ;
        RECT 56.255 161.045 56.450 161.375 ;
        RECT 56.675 161.045 56.930 161.375 ;
        RECT 56.255 160.075 56.425 161.045 ;
        RECT 57.100 160.875 57.270 161.545 ;
        RECT 57.905 161.515 59.575 162.285 ;
        RECT 59.835 161.735 60.005 162.115 ;
        RECT 60.185 161.905 60.515 162.285 ;
        RECT 59.835 161.565 60.500 161.735 ;
        RECT 60.695 161.610 60.955 162.115 ;
        RECT 54.395 159.905 56.425 160.075 ;
        RECT 56.595 159.735 56.765 160.875 ;
        RECT 56.935 159.905 57.270 160.875 ;
        RECT 57.905 160.825 58.655 161.345 ;
        RECT 58.825 160.995 59.575 161.515 ;
        RECT 59.765 161.015 60.095 161.385 ;
        RECT 60.330 161.310 60.500 161.565 ;
        RECT 60.330 160.980 60.615 161.310 ;
        RECT 60.330 160.835 60.500 160.980 ;
        RECT 57.905 159.735 59.575 160.825 ;
        RECT 59.835 160.665 60.500 160.835 ;
        RECT 60.785 160.810 60.955 161.610 ;
        RECT 61.125 161.515 62.795 162.285 ;
        RECT 62.965 161.560 63.255 162.285 ;
        RECT 63.425 161.535 64.635 162.285 ;
        RECT 59.835 159.905 60.005 160.665 ;
        RECT 60.185 159.735 60.515 160.495 ;
        RECT 60.685 159.905 60.955 160.810 ;
        RECT 61.125 160.825 61.875 161.345 ;
        RECT 62.045 160.995 62.795 161.515 ;
        RECT 61.125 159.735 62.795 160.825 ;
        RECT 62.965 159.735 63.255 160.900 ;
        RECT 63.425 160.825 63.945 161.365 ;
        RECT 64.115 160.995 64.635 161.535 ;
        RECT 64.810 161.445 65.070 162.285 ;
        RECT 65.245 161.540 65.500 162.115 ;
        RECT 65.670 161.905 66.000 162.285 ;
        RECT 66.215 161.735 66.385 162.115 ;
        RECT 65.670 161.565 66.385 161.735 ;
        RECT 63.425 159.735 64.635 160.825 ;
        RECT 64.810 159.735 65.070 160.885 ;
        RECT 65.245 160.810 65.415 161.540 ;
        RECT 65.670 161.375 65.840 161.565 ;
        RECT 66.650 161.445 66.910 162.285 ;
        RECT 67.085 161.540 67.340 162.115 ;
        RECT 67.510 161.905 67.840 162.285 ;
        RECT 68.055 161.735 68.225 162.115 ;
        RECT 67.510 161.565 68.225 161.735 ;
        RECT 68.575 161.735 68.745 162.115 ;
        RECT 68.960 161.905 69.290 162.285 ;
        RECT 68.575 161.565 69.290 161.735 ;
        RECT 65.585 161.045 65.840 161.375 ;
        RECT 65.670 160.835 65.840 161.045 ;
        RECT 66.120 161.015 66.475 161.385 ;
        RECT 65.245 159.905 65.500 160.810 ;
        RECT 65.670 160.665 66.385 160.835 ;
        RECT 65.670 159.735 66.000 160.495 ;
        RECT 66.215 159.905 66.385 160.665 ;
        RECT 66.650 159.735 66.910 160.885 ;
        RECT 67.085 160.810 67.255 161.540 ;
        RECT 67.510 161.375 67.680 161.565 ;
        RECT 67.425 161.045 67.680 161.375 ;
        RECT 67.510 160.835 67.680 161.045 ;
        RECT 67.960 161.015 68.315 161.385 ;
        RECT 68.485 161.015 68.840 161.385 ;
        RECT 69.120 161.375 69.290 161.565 ;
        RECT 69.460 161.540 69.715 162.115 ;
        RECT 69.120 161.045 69.375 161.375 ;
        RECT 69.120 160.835 69.290 161.045 ;
        RECT 67.085 159.905 67.340 160.810 ;
        RECT 67.510 160.665 68.225 160.835 ;
        RECT 67.510 159.735 67.840 160.495 ;
        RECT 68.055 159.905 68.225 160.665 ;
        RECT 68.575 160.665 69.290 160.835 ;
        RECT 69.545 160.810 69.715 161.540 ;
        RECT 69.890 161.445 70.150 162.285 ;
        RECT 70.415 161.735 70.585 162.115 ;
        RECT 70.800 161.905 71.130 162.285 ;
        RECT 70.415 161.565 71.130 161.735 ;
        RECT 70.325 161.015 70.680 161.385 ;
        RECT 70.960 161.375 71.130 161.565 ;
        RECT 71.300 161.540 71.555 162.115 ;
        RECT 70.960 161.045 71.215 161.375 ;
        RECT 68.575 159.905 68.745 160.665 ;
        RECT 68.960 159.735 69.290 160.495 ;
        RECT 69.460 159.905 69.715 160.810 ;
        RECT 69.890 159.735 70.150 160.885 ;
        RECT 70.960 160.835 71.130 161.045 ;
        RECT 70.415 160.665 71.130 160.835 ;
        RECT 71.385 160.810 71.555 161.540 ;
        RECT 71.730 161.445 71.990 162.285 ;
        RECT 72.625 161.515 75.215 162.285 ;
        RECT 75.390 161.740 80.735 162.285 ;
        RECT 70.415 159.905 70.585 160.665 ;
        RECT 70.800 159.735 71.130 160.495 ;
        RECT 71.300 159.905 71.555 160.810 ;
        RECT 71.730 159.735 71.990 160.885 ;
        RECT 72.625 160.825 73.835 161.345 ;
        RECT 74.005 160.995 75.215 161.515 ;
        RECT 72.625 159.735 75.215 160.825 ;
        RECT 76.980 160.170 77.330 161.420 ;
        RECT 78.810 160.910 79.150 161.740 ;
        RECT 80.965 161.465 81.175 162.285 ;
        RECT 81.345 161.485 81.675 162.115 ;
        RECT 81.345 160.885 81.595 161.485 ;
        RECT 81.845 161.465 82.075 162.285 ;
        RECT 82.560 161.475 82.805 162.080 ;
        RECT 83.025 161.750 83.535 162.285 ;
        RECT 82.285 161.305 83.515 161.475 ;
        RECT 81.765 161.045 82.095 161.295 ;
        RECT 75.390 159.735 80.735 160.170 ;
        RECT 80.965 159.735 81.175 160.875 ;
        RECT 81.345 159.905 81.675 160.885 ;
        RECT 81.845 159.735 82.075 160.875 ;
        RECT 82.285 160.495 82.625 161.305 ;
        RECT 82.795 160.740 83.545 160.930 ;
        RECT 82.285 160.085 82.800 160.495 ;
        RECT 83.035 159.735 83.205 160.495 ;
        RECT 83.375 160.075 83.545 160.740 ;
        RECT 83.715 160.755 83.905 162.115 ;
        RECT 84.075 161.605 84.350 162.115 ;
        RECT 84.540 161.750 85.070 162.115 ;
        RECT 85.495 161.885 85.825 162.285 ;
        RECT 84.895 161.715 85.070 161.750 ;
        RECT 84.075 161.435 84.355 161.605 ;
        RECT 84.075 160.955 84.350 161.435 ;
        RECT 84.555 160.755 84.725 161.555 ;
        RECT 83.715 160.585 84.725 160.755 ;
        RECT 84.895 161.545 85.825 161.715 ;
        RECT 85.995 161.545 86.250 162.115 ;
        RECT 86.515 161.735 86.685 162.115 ;
        RECT 86.865 161.905 87.195 162.285 ;
        RECT 86.515 161.565 87.180 161.735 ;
        RECT 87.375 161.610 87.635 162.115 ;
        RECT 84.895 160.415 85.065 161.545 ;
        RECT 85.655 161.375 85.825 161.545 ;
        RECT 83.940 160.245 85.065 160.415 ;
        RECT 85.235 161.045 85.430 161.375 ;
        RECT 85.655 161.045 85.910 161.375 ;
        RECT 85.235 160.075 85.405 161.045 ;
        RECT 86.080 160.875 86.250 161.545 ;
        RECT 86.445 161.015 86.775 161.385 ;
        RECT 87.010 161.310 87.180 161.565 ;
        RECT 83.375 159.905 85.405 160.075 ;
        RECT 85.575 159.735 85.745 160.875 ;
        RECT 85.915 159.905 86.250 160.875 ;
        RECT 87.010 160.980 87.295 161.310 ;
        RECT 87.010 160.835 87.180 160.980 ;
        RECT 86.515 160.665 87.180 160.835 ;
        RECT 87.465 160.810 87.635 161.610 ;
        RECT 88.725 161.560 89.015 162.285 ;
        RECT 90.020 161.945 90.275 162.105 ;
        RECT 89.935 161.775 90.275 161.945 ;
        RECT 90.455 161.825 90.740 162.285 ;
        RECT 90.020 161.575 90.275 161.775 ;
        RECT 86.515 159.905 86.685 160.665 ;
        RECT 86.865 159.735 87.195 160.495 ;
        RECT 87.365 159.905 87.635 160.810 ;
        RECT 88.725 159.735 89.015 160.900 ;
        RECT 90.020 160.715 90.200 161.575 ;
        RECT 90.920 161.375 91.170 162.025 ;
        RECT 90.370 161.045 91.170 161.375 ;
        RECT 90.020 160.045 90.275 160.715 ;
        RECT 90.455 159.735 90.740 160.535 ;
        RECT 90.920 160.455 91.170 161.045 ;
        RECT 91.370 161.690 91.690 162.020 ;
        RECT 91.870 161.805 92.530 162.285 ;
        RECT 92.730 161.895 93.580 162.065 ;
        RECT 91.370 160.795 91.560 161.690 ;
        RECT 91.880 161.365 92.540 161.635 ;
        RECT 92.210 161.305 92.540 161.365 ;
        RECT 91.730 161.135 92.060 161.195 ;
        RECT 92.730 161.135 92.900 161.895 ;
        RECT 94.140 161.825 94.460 162.285 ;
        RECT 94.660 161.645 94.910 162.075 ;
        RECT 95.200 161.845 95.610 162.285 ;
        RECT 95.780 161.905 96.795 162.105 ;
        RECT 93.070 161.475 94.320 161.645 ;
        RECT 93.070 161.355 93.400 161.475 ;
        RECT 91.730 160.965 93.630 161.135 ;
        RECT 91.370 160.625 93.290 160.795 ;
        RECT 91.370 160.605 91.690 160.625 ;
        RECT 90.920 159.945 91.250 160.455 ;
        RECT 91.520 159.995 91.690 160.605 ;
        RECT 93.460 160.455 93.630 160.965 ;
        RECT 93.800 160.895 93.980 161.305 ;
        RECT 94.150 160.715 94.320 161.475 ;
        RECT 91.860 159.735 92.190 160.425 ;
        RECT 92.420 160.285 93.630 160.455 ;
        RECT 93.800 160.405 94.320 160.715 ;
        RECT 94.490 161.305 94.910 161.645 ;
        RECT 95.200 161.305 95.610 161.635 ;
        RECT 94.490 160.535 94.680 161.305 ;
        RECT 95.780 161.175 95.950 161.905 ;
        RECT 97.095 161.735 97.265 162.065 ;
        RECT 97.435 161.905 97.765 162.285 ;
        RECT 96.120 161.355 96.470 161.725 ;
        RECT 95.780 161.135 96.200 161.175 ;
        RECT 94.850 160.965 96.200 161.135 ;
        RECT 94.850 160.805 95.100 160.965 ;
        RECT 95.610 160.535 95.860 160.795 ;
        RECT 94.490 160.285 95.860 160.535 ;
        RECT 92.420 159.995 92.660 160.285 ;
        RECT 93.460 160.205 93.630 160.285 ;
        RECT 92.860 159.735 93.280 160.115 ;
        RECT 93.460 159.955 94.090 160.205 ;
        RECT 94.560 159.735 94.890 160.115 ;
        RECT 95.060 159.995 95.230 160.285 ;
        RECT 96.030 160.120 96.200 160.965 ;
        RECT 96.650 160.795 96.870 161.665 ;
        RECT 97.095 161.545 97.790 161.735 ;
        RECT 96.370 160.415 96.870 160.795 ;
        RECT 97.040 160.745 97.450 161.365 ;
        RECT 97.620 160.575 97.790 161.545 ;
        RECT 97.095 160.405 97.790 160.575 ;
        RECT 95.410 159.735 95.790 160.115 ;
        RECT 96.030 159.950 96.860 160.120 ;
        RECT 97.095 159.905 97.265 160.405 ;
        RECT 97.435 159.735 97.765 160.235 ;
        RECT 97.980 159.905 98.205 162.025 ;
        RECT 98.375 161.905 98.705 162.285 ;
        RECT 98.875 161.735 99.045 162.025 ;
        RECT 99.405 161.820 99.655 162.285 ;
        RECT 98.380 161.565 99.045 161.735 ;
        RECT 99.825 161.645 99.995 162.115 ;
        RECT 100.245 161.825 100.415 162.285 ;
        RECT 100.665 161.645 100.835 162.115 ;
        RECT 101.085 161.825 101.255 162.285 ;
        RECT 101.505 161.645 101.675 162.115 ;
        RECT 102.045 161.825 102.310 162.285 ;
        RECT 98.380 160.575 98.610 161.565 ;
        RECT 99.305 161.465 101.675 161.645 ;
        RECT 102.640 161.655 102.925 162.115 ;
        RECT 103.095 161.825 103.365 162.285 ;
        RECT 102.640 161.485 103.595 161.655 ;
        RECT 98.780 160.745 99.130 161.395 ;
        RECT 99.305 160.875 99.655 161.465 ;
        RECT 99.825 161.045 102.335 161.295 ;
        RECT 99.305 160.705 101.755 160.875 ;
        RECT 99.305 160.685 100.075 160.705 ;
        RECT 98.380 160.405 99.045 160.575 ;
        RECT 98.375 159.735 98.705 160.235 ;
        RECT 98.875 159.905 99.045 160.405 ;
        RECT 99.405 159.735 99.575 160.195 ;
        RECT 99.745 159.905 100.075 160.685 ;
        RECT 100.245 159.735 100.415 160.535 ;
        RECT 100.585 159.905 100.915 160.705 ;
        RECT 101.085 159.735 101.255 160.535 ;
        RECT 101.425 159.905 101.755 160.705 ;
        RECT 102.015 159.735 102.310 160.875 ;
        RECT 102.525 160.755 103.215 161.315 ;
        RECT 103.385 160.585 103.595 161.485 ;
        RECT 102.640 160.365 103.595 160.585 ;
        RECT 103.765 161.315 104.165 162.115 ;
        RECT 104.355 161.655 104.635 162.115 ;
        RECT 105.155 161.825 105.480 162.285 ;
        RECT 104.355 161.485 105.480 161.655 ;
        RECT 105.650 161.545 106.035 162.115 ;
        RECT 105.030 161.375 105.480 161.485 ;
        RECT 103.765 160.755 104.860 161.315 ;
        RECT 105.030 161.045 105.585 161.375 ;
        RECT 102.640 159.905 102.925 160.365 ;
        RECT 103.095 159.735 103.365 160.195 ;
        RECT 103.765 159.905 104.165 160.755 ;
        RECT 105.030 160.585 105.480 161.045 ;
        RECT 105.755 160.875 106.035 161.545 ;
        RECT 106.780 161.655 107.065 162.115 ;
        RECT 107.235 161.825 107.505 162.285 ;
        RECT 106.780 161.485 107.735 161.655 ;
        RECT 104.355 160.365 105.480 160.585 ;
        RECT 104.355 159.905 104.635 160.365 ;
        RECT 105.155 159.735 105.480 160.195 ;
        RECT 105.650 159.905 106.035 160.875 ;
        RECT 106.665 160.755 107.355 161.315 ;
        RECT 107.525 160.585 107.735 161.485 ;
        RECT 106.780 160.365 107.735 160.585 ;
        RECT 107.905 161.315 108.305 162.115 ;
        RECT 108.495 161.655 108.775 162.115 ;
        RECT 109.295 161.825 109.620 162.285 ;
        RECT 108.495 161.485 109.620 161.655 ;
        RECT 109.790 161.545 110.175 162.115 ;
        RECT 109.170 161.375 109.620 161.485 ;
        RECT 107.905 160.755 109.000 161.315 ;
        RECT 109.170 161.045 109.725 161.375 ;
        RECT 106.780 159.905 107.065 160.365 ;
        RECT 107.235 159.735 107.505 160.195 ;
        RECT 107.905 159.905 108.305 160.755 ;
        RECT 109.170 160.585 109.620 161.045 ;
        RECT 109.895 160.875 110.175 161.545 ;
        RECT 110.620 161.475 110.865 162.080 ;
        RECT 111.085 161.750 111.595 162.285 ;
        RECT 108.495 160.365 109.620 160.585 ;
        RECT 108.495 159.905 108.775 160.365 ;
        RECT 109.295 159.735 109.620 160.195 ;
        RECT 109.790 159.905 110.175 160.875 ;
        RECT 110.345 161.305 111.575 161.475 ;
        RECT 110.345 160.495 110.685 161.305 ;
        RECT 110.855 160.740 111.605 160.930 ;
        RECT 110.345 160.085 110.860 160.495 ;
        RECT 111.095 159.735 111.265 160.495 ;
        RECT 111.435 160.075 111.605 160.740 ;
        RECT 111.775 160.755 111.965 162.115 ;
        RECT 112.135 161.265 112.410 162.115 ;
        RECT 112.600 161.750 113.130 162.115 ;
        RECT 113.555 161.885 113.885 162.285 ;
        RECT 112.955 161.715 113.130 161.750 ;
        RECT 112.135 161.095 112.415 161.265 ;
        RECT 112.135 160.955 112.410 161.095 ;
        RECT 112.615 160.755 112.785 161.555 ;
        RECT 111.775 160.585 112.785 160.755 ;
        RECT 112.955 161.545 113.885 161.715 ;
        RECT 114.055 161.545 114.310 162.115 ;
        RECT 114.485 161.560 114.775 162.285 ;
        RECT 112.955 160.415 113.125 161.545 ;
        RECT 113.715 161.375 113.885 161.545 ;
        RECT 112.000 160.245 113.125 160.415 ;
        RECT 113.295 161.045 113.490 161.375 ;
        RECT 113.715 161.045 113.970 161.375 ;
        RECT 113.295 160.075 113.465 161.045 ;
        RECT 114.140 160.875 114.310 161.545 ;
        RECT 115.220 161.475 115.465 162.080 ;
        RECT 115.685 161.750 116.195 162.285 ;
        RECT 114.945 161.305 116.175 161.475 ;
        RECT 111.435 159.905 113.465 160.075 ;
        RECT 113.635 159.735 113.805 160.875 ;
        RECT 113.975 159.905 114.310 160.875 ;
        RECT 114.485 159.735 114.775 160.900 ;
        RECT 114.945 160.495 115.285 161.305 ;
        RECT 115.455 160.740 116.205 160.930 ;
        RECT 114.945 160.085 115.460 160.495 ;
        RECT 115.695 159.735 115.865 160.495 ;
        RECT 116.035 160.075 116.205 160.740 ;
        RECT 116.375 160.755 116.565 162.115 ;
        RECT 116.735 161.945 117.010 162.115 ;
        RECT 116.735 161.775 117.015 161.945 ;
        RECT 116.735 160.955 117.010 161.775 ;
        RECT 117.200 161.750 117.730 162.115 ;
        RECT 118.155 161.885 118.485 162.285 ;
        RECT 117.555 161.715 117.730 161.750 ;
        RECT 117.215 160.755 117.385 161.555 ;
        RECT 116.375 160.585 117.385 160.755 ;
        RECT 117.555 161.545 118.485 161.715 ;
        RECT 118.655 161.545 118.910 162.115 ;
        RECT 117.555 160.415 117.725 161.545 ;
        RECT 118.315 161.375 118.485 161.545 ;
        RECT 116.600 160.245 117.725 160.415 ;
        RECT 117.895 161.045 118.090 161.375 ;
        RECT 118.315 161.045 118.570 161.375 ;
        RECT 117.895 160.075 118.065 161.045 ;
        RECT 118.740 160.875 118.910 161.545 ;
        RECT 119.125 161.465 119.355 162.285 ;
        RECT 119.525 161.485 119.855 162.115 ;
        RECT 119.105 161.045 119.435 161.295 ;
        RECT 119.605 160.885 119.855 161.485 ;
        RECT 120.025 161.465 120.235 162.285 ;
        RECT 121.015 161.735 121.185 162.115 ;
        RECT 121.365 161.905 121.695 162.285 ;
        RECT 121.015 161.565 121.680 161.735 ;
        RECT 121.875 161.610 122.135 162.115 ;
        RECT 120.945 161.015 121.275 161.385 ;
        RECT 121.510 161.310 121.680 161.565 ;
        RECT 116.035 159.905 118.065 160.075 ;
        RECT 118.235 159.735 118.405 160.875 ;
        RECT 118.575 159.905 118.910 160.875 ;
        RECT 119.125 159.735 119.355 160.875 ;
        RECT 119.525 159.905 119.855 160.885 ;
        RECT 121.510 160.980 121.795 161.310 ;
        RECT 120.025 159.735 120.235 160.875 ;
        RECT 121.510 160.835 121.680 160.980 ;
        RECT 121.015 160.665 121.680 160.835 ;
        RECT 121.965 160.810 122.135 161.610 ;
        RECT 122.765 161.515 126.275 162.285 ;
        RECT 126.445 161.535 127.655 162.285 ;
        RECT 121.015 159.905 121.185 160.665 ;
        RECT 121.365 159.735 121.695 160.495 ;
        RECT 121.865 159.905 122.135 160.810 ;
        RECT 122.765 160.825 124.455 161.345 ;
        RECT 124.625 160.995 126.275 161.515 ;
        RECT 126.445 160.825 126.965 161.365 ;
        RECT 127.135 160.995 127.655 161.535 ;
        RECT 122.765 159.735 126.275 160.825 ;
        RECT 126.445 159.735 127.655 160.825 ;
        RECT 14.580 159.565 127.740 159.735 ;
        RECT 14.665 158.475 15.875 159.565 ;
        RECT 14.665 157.765 15.185 158.305 ;
        RECT 15.355 157.935 15.875 158.475 ;
        RECT 16.045 158.475 17.255 159.565 ;
        RECT 16.045 157.935 16.565 158.475 ;
        RECT 17.485 158.425 17.695 159.565 ;
        RECT 17.865 158.415 18.195 159.395 ;
        RECT 18.365 158.425 18.595 159.565 ;
        RECT 18.845 158.425 19.075 159.565 ;
        RECT 19.245 158.415 19.575 159.395 ;
        RECT 19.745 158.425 19.955 159.565 ;
        RECT 20.185 158.805 20.700 159.215 ;
        RECT 20.935 158.805 21.105 159.565 ;
        RECT 21.275 159.225 23.305 159.395 ;
        RECT 16.735 157.765 17.255 158.305 ;
        RECT 14.665 157.015 15.875 157.765 ;
        RECT 16.045 157.015 17.255 157.765 ;
        RECT 17.485 157.015 17.695 157.835 ;
        RECT 17.865 157.815 18.115 158.415 ;
        RECT 18.285 158.005 18.615 158.255 ;
        RECT 18.825 158.005 19.155 158.255 ;
        RECT 17.865 157.185 18.195 157.815 ;
        RECT 18.365 157.015 18.595 157.835 ;
        RECT 18.845 157.015 19.075 157.835 ;
        RECT 19.325 157.815 19.575 158.415 ;
        RECT 20.185 157.995 20.525 158.805 ;
        RECT 21.275 158.560 21.445 159.225 ;
        RECT 21.840 158.885 22.965 159.055 ;
        RECT 20.695 158.370 21.445 158.560 ;
        RECT 21.615 158.545 22.625 158.715 ;
        RECT 19.245 157.185 19.575 157.815 ;
        RECT 19.745 157.015 19.955 157.835 ;
        RECT 20.185 157.825 21.415 157.995 ;
        RECT 20.460 157.220 20.705 157.825 ;
        RECT 20.925 157.015 21.435 157.550 ;
        RECT 21.615 157.185 21.805 158.545 ;
        RECT 21.975 157.525 22.250 158.345 ;
        RECT 22.455 157.745 22.625 158.545 ;
        RECT 22.795 157.755 22.965 158.885 ;
        RECT 23.135 158.255 23.305 159.225 ;
        RECT 23.475 158.425 23.645 159.565 ;
        RECT 23.815 158.425 24.150 159.395 ;
        RECT 23.135 157.925 23.330 158.255 ;
        RECT 23.555 157.925 23.810 158.255 ;
        RECT 23.555 157.755 23.725 157.925 ;
        RECT 23.980 157.755 24.150 158.425 ;
        RECT 24.325 158.400 24.615 159.565 ;
        RECT 24.875 158.635 25.045 159.395 ;
        RECT 25.225 158.805 25.555 159.565 ;
        RECT 24.875 158.465 25.540 158.635 ;
        RECT 25.725 158.490 25.995 159.395 ;
        RECT 25.370 158.320 25.540 158.465 ;
        RECT 24.805 157.915 25.135 158.285 ;
        RECT 25.370 157.990 25.655 158.320 ;
        RECT 22.795 157.585 23.725 157.755 ;
        RECT 22.795 157.550 22.970 157.585 ;
        RECT 21.975 157.355 22.255 157.525 ;
        RECT 21.975 157.185 22.250 157.355 ;
        RECT 22.440 157.185 22.970 157.550 ;
        RECT 23.395 157.015 23.725 157.415 ;
        RECT 23.895 157.185 24.150 157.755 ;
        RECT 24.325 157.015 24.615 157.740 ;
        RECT 25.370 157.735 25.540 157.990 ;
        RECT 24.875 157.565 25.540 157.735 ;
        RECT 25.825 157.690 25.995 158.490 ;
        RECT 26.165 158.475 27.835 159.565 ;
        RECT 28.120 158.935 28.405 159.395 ;
        RECT 28.575 159.105 28.845 159.565 ;
        RECT 28.120 158.715 29.075 158.935 ;
        RECT 26.165 157.955 26.915 158.475 ;
        RECT 27.085 157.785 27.835 158.305 ;
        RECT 28.005 157.985 28.695 158.545 ;
        RECT 28.865 157.815 29.075 158.715 ;
        RECT 24.875 157.185 25.045 157.565 ;
        RECT 25.225 157.015 25.555 157.395 ;
        RECT 25.735 157.185 25.995 157.690 ;
        RECT 26.165 157.015 27.835 157.785 ;
        RECT 28.120 157.645 29.075 157.815 ;
        RECT 29.245 158.545 29.645 159.395 ;
        RECT 29.835 158.935 30.115 159.395 ;
        RECT 30.635 159.105 30.960 159.565 ;
        RECT 29.835 158.715 30.960 158.935 ;
        RECT 29.245 157.985 30.340 158.545 ;
        RECT 30.510 158.255 30.960 158.715 ;
        RECT 31.130 158.425 31.515 159.395 ;
        RECT 31.800 158.935 32.085 159.395 ;
        RECT 32.255 159.105 32.525 159.565 ;
        RECT 31.800 158.715 32.755 158.935 ;
        RECT 28.120 157.185 28.405 157.645 ;
        RECT 28.575 157.015 28.845 157.475 ;
        RECT 29.245 157.185 29.645 157.985 ;
        RECT 30.510 157.925 31.065 158.255 ;
        RECT 30.510 157.815 30.960 157.925 ;
        RECT 29.835 157.645 30.960 157.815 ;
        RECT 31.235 157.755 31.515 158.425 ;
        RECT 31.685 157.985 32.375 158.545 ;
        RECT 32.545 157.815 32.755 158.715 ;
        RECT 29.835 157.185 30.115 157.645 ;
        RECT 30.635 157.015 30.960 157.475 ;
        RECT 31.130 157.185 31.515 157.755 ;
        RECT 31.800 157.645 32.755 157.815 ;
        RECT 32.925 158.545 33.325 159.395 ;
        RECT 33.515 158.935 33.795 159.395 ;
        RECT 34.315 159.105 34.640 159.565 ;
        RECT 33.515 158.715 34.640 158.935 ;
        RECT 32.925 157.985 34.020 158.545 ;
        RECT 34.190 158.255 34.640 158.715 ;
        RECT 34.810 158.425 35.195 159.395 ;
        RECT 31.800 157.185 32.085 157.645 ;
        RECT 32.255 157.015 32.525 157.475 ;
        RECT 32.925 157.185 33.325 157.985 ;
        RECT 34.190 157.925 34.745 158.255 ;
        RECT 34.190 157.815 34.640 157.925 ;
        RECT 33.515 157.645 34.640 157.815 ;
        RECT 34.915 157.755 35.195 158.425 ;
        RECT 35.365 158.475 38.875 159.565 ;
        RECT 39.250 158.595 39.580 159.395 ;
        RECT 39.750 158.765 40.080 159.565 ;
        RECT 40.380 158.595 40.710 159.395 ;
        RECT 41.355 158.765 41.605 159.565 ;
        RECT 35.365 157.955 37.055 158.475 ;
        RECT 39.250 158.425 41.685 158.595 ;
        RECT 41.875 158.425 42.045 159.565 ;
        RECT 42.215 158.425 42.555 159.395 ;
        RECT 42.930 158.595 43.260 159.395 ;
        RECT 43.430 158.765 43.760 159.565 ;
        RECT 44.060 158.595 44.390 159.395 ;
        RECT 45.035 158.765 45.285 159.565 ;
        RECT 42.930 158.425 45.365 158.595 ;
        RECT 45.555 158.425 45.725 159.565 ;
        RECT 45.895 158.425 46.235 159.395 ;
        RECT 46.520 158.935 46.805 159.395 ;
        RECT 46.975 159.105 47.245 159.565 ;
        RECT 46.520 158.715 47.475 158.935 ;
        RECT 37.225 157.785 38.875 158.305 ;
        RECT 39.045 158.005 39.395 158.255 ;
        RECT 39.580 157.795 39.750 158.425 ;
        RECT 39.920 158.005 40.250 158.205 ;
        RECT 40.420 158.005 40.750 158.205 ;
        RECT 40.920 158.005 41.340 158.205 ;
        RECT 41.515 158.175 41.685 158.425 ;
        RECT 41.515 158.005 42.210 158.175 ;
        RECT 33.515 157.185 33.795 157.645 ;
        RECT 34.315 157.015 34.640 157.475 ;
        RECT 34.810 157.185 35.195 157.755 ;
        RECT 35.365 157.015 38.875 157.785 ;
        RECT 39.250 157.185 39.750 157.795 ;
        RECT 40.380 157.665 41.605 157.835 ;
        RECT 42.380 157.815 42.555 158.425 ;
        RECT 42.725 158.005 43.075 158.255 ;
        RECT 40.380 157.185 40.710 157.665 ;
        RECT 40.880 157.015 41.105 157.475 ;
        RECT 41.275 157.185 41.605 157.665 ;
        RECT 41.795 157.015 42.045 157.815 ;
        RECT 42.215 157.185 42.555 157.815 ;
        RECT 43.260 157.795 43.430 158.425 ;
        RECT 43.600 158.005 43.930 158.205 ;
        RECT 44.100 158.005 44.430 158.205 ;
        RECT 44.600 158.005 45.020 158.205 ;
        RECT 45.195 158.175 45.365 158.425 ;
        RECT 45.195 158.005 45.890 158.175 ;
        RECT 42.930 157.185 43.430 157.795 ;
        RECT 44.060 157.665 45.285 157.835 ;
        RECT 46.060 157.815 46.235 158.425 ;
        RECT 46.405 157.985 47.095 158.545 ;
        RECT 47.265 157.815 47.475 158.715 ;
        RECT 44.060 157.185 44.390 157.665 ;
        RECT 44.560 157.015 44.785 157.475 ;
        RECT 44.955 157.185 45.285 157.665 ;
        RECT 45.475 157.015 45.725 157.815 ;
        RECT 45.895 157.185 46.235 157.815 ;
        RECT 46.520 157.645 47.475 157.815 ;
        RECT 47.645 158.545 48.045 159.395 ;
        RECT 48.235 158.935 48.515 159.395 ;
        RECT 49.035 159.105 49.360 159.565 ;
        RECT 48.235 158.715 49.360 158.935 ;
        RECT 47.645 157.985 48.740 158.545 ;
        RECT 48.910 158.255 49.360 158.715 ;
        RECT 49.530 158.425 49.915 159.395 ;
        RECT 46.520 157.185 46.805 157.645 ;
        RECT 46.975 157.015 47.245 157.475 ;
        RECT 47.645 157.185 48.045 157.985 ;
        RECT 48.910 157.925 49.465 158.255 ;
        RECT 48.910 157.815 49.360 157.925 ;
        RECT 48.235 157.645 49.360 157.815 ;
        RECT 49.635 157.755 49.915 158.425 ;
        RECT 50.085 158.400 50.375 159.565 ;
        RECT 50.545 158.425 50.885 159.395 ;
        RECT 51.055 158.425 51.225 159.565 ;
        RECT 51.495 158.765 51.745 159.565 ;
        RECT 52.390 158.595 52.720 159.395 ;
        RECT 53.020 158.765 53.350 159.565 ;
        RECT 53.520 158.595 53.850 159.395 ;
        RECT 54.690 159.130 60.035 159.565 ;
        RECT 51.415 158.425 53.850 158.595 ;
        RECT 48.235 157.185 48.515 157.645 ;
        RECT 49.035 157.015 49.360 157.475 ;
        RECT 49.530 157.185 49.915 157.755 ;
        RECT 50.545 157.815 50.720 158.425 ;
        RECT 51.415 158.175 51.585 158.425 ;
        RECT 50.890 158.005 51.585 158.175 ;
        RECT 51.760 158.005 52.180 158.205 ;
        RECT 52.350 158.005 52.680 158.205 ;
        RECT 52.850 158.005 53.180 158.205 ;
        RECT 50.085 157.015 50.375 157.740 ;
        RECT 50.545 157.185 50.885 157.815 ;
        RECT 51.055 157.015 51.305 157.815 ;
        RECT 51.495 157.665 52.720 157.835 ;
        RECT 51.495 157.185 51.825 157.665 ;
        RECT 51.995 157.015 52.220 157.475 ;
        RECT 52.390 157.185 52.720 157.665 ;
        RECT 53.350 157.795 53.520 158.425 ;
        RECT 53.705 158.005 54.055 158.255 ;
        RECT 56.280 157.880 56.630 159.130 ;
        RECT 60.265 158.425 60.475 159.565 ;
        RECT 60.645 158.415 60.975 159.395 ;
        RECT 61.145 158.425 61.375 159.565 ;
        RECT 61.735 158.415 62.065 159.565 ;
        RECT 62.235 158.545 62.405 159.395 ;
        RECT 62.575 158.765 62.905 159.565 ;
        RECT 63.075 158.545 63.245 159.395 ;
        RECT 63.425 158.765 63.665 159.565 ;
        RECT 63.835 158.585 64.165 159.395 ;
        RECT 53.350 157.185 53.850 157.795 ;
        RECT 58.110 157.560 58.450 158.390 ;
        RECT 54.690 157.015 60.035 157.560 ;
        RECT 60.265 157.015 60.475 157.835 ;
        RECT 60.645 157.815 60.895 158.415 ;
        RECT 62.235 158.375 63.245 158.545 ;
        RECT 63.450 158.415 64.165 158.585 ;
        RECT 64.805 158.475 68.315 159.565 ;
        RECT 68.575 158.635 68.745 159.395 ;
        RECT 68.960 158.805 69.290 159.565 ;
        RECT 61.065 158.005 61.395 158.255 ;
        RECT 62.235 158.205 62.730 158.375 ;
        RECT 62.235 158.035 62.735 158.205 ;
        RECT 63.450 158.175 63.620 158.415 ;
        RECT 62.235 157.835 62.730 158.035 ;
        RECT 63.120 158.005 63.620 158.175 ;
        RECT 63.790 158.005 64.170 158.245 ;
        RECT 63.450 157.835 63.620 158.005 ;
        RECT 64.805 157.955 66.495 158.475 ;
        RECT 68.575 158.465 69.290 158.635 ;
        RECT 69.460 158.490 69.715 159.395 ;
        RECT 60.645 157.185 60.975 157.815 ;
        RECT 61.145 157.015 61.375 157.835 ;
        RECT 61.735 157.015 62.065 157.815 ;
        RECT 62.235 157.665 63.245 157.835 ;
        RECT 63.450 157.665 64.085 157.835 ;
        RECT 66.665 157.785 68.315 158.305 ;
        RECT 68.485 157.915 68.840 158.285 ;
        RECT 69.120 158.255 69.290 158.465 ;
        RECT 69.120 157.925 69.375 158.255 ;
        RECT 62.235 157.185 62.405 157.665 ;
        RECT 62.575 157.015 62.905 157.495 ;
        RECT 63.075 157.185 63.245 157.665 ;
        RECT 63.495 157.015 63.735 157.495 ;
        RECT 63.915 157.185 64.085 157.665 ;
        RECT 64.805 157.015 68.315 157.785 ;
        RECT 69.120 157.735 69.290 157.925 ;
        RECT 69.545 157.760 69.715 158.490 ;
        RECT 69.890 158.415 70.150 159.565 ;
        RECT 70.415 158.635 70.585 159.395 ;
        RECT 70.800 158.805 71.130 159.565 ;
        RECT 70.415 158.465 71.130 158.635 ;
        RECT 71.300 158.490 71.555 159.395 ;
        RECT 70.325 157.915 70.680 158.285 ;
        RECT 70.960 158.255 71.130 158.465 ;
        RECT 70.960 157.925 71.215 158.255 ;
        RECT 68.575 157.565 69.290 157.735 ;
        RECT 68.575 157.185 68.745 157.565 ;
        RECT 68.960 157.015 69.290 157.395 ;
        RECT 69.460 157.185 69.715 157.760 ;
        RECT 69.890 157.015 70.150 157.855 ;
        RECT 70.960 157.735 71.130 157.925 ;
        RECT 71.385 157.760 71.555 158.490 ;
        RECT 71.730 158.415 71.990 159.565 ;
        RECT 72.370 158.595 72.700 159.395 ;
        RECT 72.870 158.765 73.200 159.565 ;
        RECT 73.500 158.595 73.830 159.395 ;
        RECT 74.475 158.765 74.725 159.565 ;
        RECT 72.370 158.425 74.805 158.595 ;
        RECT 74.995 158.425 75.165 159.565 ;
        RECT 75.335 158.425 75.675 159.395 ;
        RECT 72.165 158.005 72.515 158.255 ;
        RECT 70.415 157.565 71.130 157.735 ;
        RECT 70.415 157.185 70.585 157.565 ;
        RECT 70.800 157.015 71.130 157.395 ;
        RECT 71.300 157.185 71.555 157.760 ;
        RECT 71.730 157.015 71.990 157.855 ;
        RECT 72.700 157.795 72.870 158.425 ;
        RECT 73.040 158.005 73.370 158.205 ;
        RECT 73.540 158.005 73.870 158.205 ;
        RECT 74.040 158.005 74.460 158.205 ;
        RECT 74.635 158.175 74.805 158.425 ;
        RECT 74.635 158.005 75.330 158.175 ;
        RECT 72.370 157.185 72.870 157.795 ;
        RECT 73.500 157.665 74.725 157.835 ;
        RECT 75.500 157.815 75.675 158.425 ;
        RECT 75.845 158.400 76.135 159.565 ;
        RECT 76.970 158.595 77.300 159.395 ;
        RECT 77.470 158.765 77.800 159.565 ;
        RECT 78.100 158.595 78.430 159.395 ;
        RECT 79.075 158.765 79.325 159.565 ;
        RECT 76.970 158.425 79.405 158.595 ;
        RECT 79.595 158.425 79.765 159.565 ;
        RECT 79.935 158.425 80.275 159.395 ;
        RECT 81.280 159.225 81.535 159.255 ;
        RECT 81.195 159.055 81.535 159.225 ;
        RECT 76.765 158.005 77.115 158.255 ;
        RECT 73.500 157.185 73.830 157.665 ;
        RECT 74.000 157.015 74.225 157.475 ;
        RECT 74.395 157.185 74.725 157.665 ;
        RECT 74.915 157.015 75.165 157.815 ;
        RECT 75.335 157.185 75.675 157.815 ;
        RECT 77.300 157.795 77.470 158.425 ;
        RECT 77.640 158.005 77.970 158.205 ;
        RECT 78.140 158.005 78.470 158.205 ;
        RECT 78.640 158.005 79.060 158.205 ;
        RECT 79.235 158.175 79.405 158.425 ;
        RECT 79.235 158.005 79.930 158.175 ;
        RECT 75.845 157.015 76.135 157.740 ;
        RECT 76.970 157.185 77.470 157.795 ;
        RECT 78.100 157.665 79.325 157.835 ;
        RECT 80.100 157.815 80.275 158.425 ;
        RECT 78.100 157.185 78.430 157.665 ;
        RECT 78.600 157.015 78.825 157.475 ;
        RECT 78.995 157.185 79.325 157.665 ;
        RECT 79.515 157.015 79.765 157.815 ;
        RECT 79.935 157.185 80.275 157.815 ;
        RECT 81.280 158.585 81.535 159.055 ;
        RECT 81.715 158.765 82.000 159.565 ;
        RECT 82.180 158.845 82.510 159.355 ;
        RECT 81.280 157.725 81.460 158.585 ;
        RECT 82.180 158.255 82.430 158.845 ;
        RECT 82.780 158.695 82.950 159.305 ;
        RECT 83.120 158.875 83.450 159.565 ;
        RECT 83.680 159.015 83.920 159.305 ;
        RECT 84.120 159.185 84.540 159.565 ;
        RECT 84.720 159.095 85.350 159.345 ;
        RECT 85.820 159.185 86.150 159.565 ;
        RECT 84.720 159.015 84.890 159.095 ;
        RECT 86.320 159.015 86.490 159.305 ;
        RECT 86.670 159.185 87.050 159.565 ;
        RECT 87.290 159.180 88.120 159.350 ;
        RECT 83.680 158.845 84.890 159.015 ;
        RECT 81.630 157.925 82.430 158.255 ;
        RECT 81.280 157.195 81.535 157.725 ;
        RECT 81.715 157.015 82.000 157.475 ;
        RECT 82.180 157.275 82.430 157.925 ;
        RECT 82.630 158.675 82.950 158.695 ;
        RECT 82.630 158.505 84.550 158.675 ;
        RECT 82.630 157.610 82.820 158.505 ;
        RECT 84.720 158.335 84.890 158.845 ;
        RECT 85.060 158.585 85.580 158.895 ;
        RECT 82.990 158.165 84.890 158.335 ;
        RECT 82.990 158.105 83.320 158.165 ;
        RECT 83.470 157.935 83.800 157.995 ;
        RECT 83.140 157.665 83.800 157.935 ;
        RECT 82.630 157.280 82.950 157.610 ;
        RECT 83.130 157.015 83.790 157.495 ;
        RECT 83.990 157.405 84.160 158.165 ;
        RECT 85.060 157.995 85.240 158.405 ;
        RECT 84.330 157.825 84.660 157.945 ;
        RECT 85.410 157.825 85.580 158.585 ;
        RECT 84.330 157.655 85.580 157.825 ;
        RECT 85.750 158.765 87.120 159.015 ;
        RECT 85.750 157.995 85.940 158.765 ;
        RECT 86.870 158.505 87.120 158.765 ;
        RECT 86.110 158.335 86.360 158.495 ;
        RECT 87.290 158.335 87.460 159.180 ;
        RECT 88.355 158.895 88.525 159.395 ;
        RECT 88.695 159.065 89.025 159.565 ;
        RECT 87.630 158.505 88.130 158.885 ;
        RECT 88.355 158.725 89.050 158.895 ;
        RECT 86.110 158.165 87.460 158.335 ;
        RECT 87.040 158.125 87.460 158.165 ;
        RECT 85.750 157.655 86.170 157.995 ;
        RECT 86.460 157.665 86.870 157.995 ;
        RECT 83.990 157.235 84.840 157.405 ;
        RECT 85.400 157.015 85.720 157.475 ;
        RECT 85.920 157.225 86.170 157.655 ;
        RECT 86.460 157.015 86.870 157.455 ;
        RECT 87.040 157.395 87.210 158.125 ;
        RECT 87.380 157.575 87.730 157.945 ;
        RECT 87.910 157.635 88.130 158.505 ;
        RECT 88.300 157.935 88.710 158.555 ;
        RECT 88.880 157.755 89.050 158.725 ;
        RECT 88.355 157.565 89.050 157.755 ;
        RECT 87.040 157.195 88.055 157.395 ;
        RECT 88.355 157.235 88.525 157.565 ;
        RECT 88.695 157.015 89.025 157.395 ;
        RECT 89.240 157.275 89.465 159.395 ;
        RECT 89.635 159.065 89.965 159.565 ;
        RECT 90.135 158.895 90.305 159.395 ;
        RECT 89.640 158.725 90.305 158.895 ;
        RECT 89.640 157.735 89.870 158.725 ;
        RECT 90.040 157.905 90.390 158.555 ;
        RECT 91.025 158.475 92.695 159.565 ;
        RECT 91.025 157.955 91.775 158.475 ;
        RECT 92.905 158.425 93.135 159.565 ;
        RECT 93.305 158.415 93.635 159.395 ;
        RECT 93.805 158.425 94.015 159.565 ;
        RECT 94.705 158.475 96.375 159.565 ;
        RECT 96.635 158.635 96.805 159.395 ;
        RECT 96.985 158.805 97.315 159.565 ;
        RECT 91.945 157.785 92.695 158.305 ;
        RECT 92.885 158.005 93.215 158.255 ;
        RECT 89.640 157.565 90.305 157.735 ;
        RECT 89.635 157.015 89.965 157.395 ;
        RECT 90.135 157.275 90.305 157.565 ;
        RECT 91.025 157.015 92.695 157.785 ;
        RECT 92.905 157.015 93.135 157.835 ;
        RECT 93.385 157.815 93.635 158.415 ;
        RECT 94.705 157.955 95.455 158.475 ;
        RECT 96.635 158.465 97.300 158.635 ;
        RECT 97.485 158.490 97.755 159.395 ;
        RECT 97.130 158.320 97.300 158.465 ;
        RECT 93.305 157.185 93.635 157.815 ;
        RECT 93.805 157.015 94.015 157.835 ;
        RECT 95.625 157.785 96.375 158.305 ;
        RECT 96.565 157.915 96.895 158.285 ;
        RECT 97.130 157.990 97.415 158.320 ;
        RECT 94.705 157.015 96.375 157.785 ;
        RECT 97.130 157.735 97.300 157.990 ;
        RECT 96.635 157.565 97.300 157.735 ;
        RECT 97.585 157.690 97.755 158.490 ;
        RECT 97.925 158.475 99.595 159.565 ;
        RECT 97.925 157.955 98.675 158.475 ;
        RECT 99.805 158.425 100.035 159.565 ;
        RECT 100.205 158.415 100.535 159.395 ;
        RECT 100.705 158.425 100.915 159.565 ;
        RECT 98.845 157.785 99.595 158.305 ;
        RECT 99.785 158.005 100.115 158.255 ;
        RECT 96.635 157.185 96.805 157.565 ;
        RECT 96.985 157.015 97.315 157.395 ;
        RECT 97.495 157.185 97.755 157.690 ;
        RECT 97.925 157.015 99.595 157.785 ;
        RECT 99.805 157.015 100.035 157.835 ;
        RECT 100.285 157.815 100.535 158.415 ;
        RECT 101.605 158.400 101.895 159.565 ;
        RECT 102.525 158.475 104.195 159.565 ;
        RECT 104.365 158.490 104.635 159.395 ;
        RECT 104.805 158.805 105.135 159.565 ;
        RECT 105.315 158.635 105.485 159.395 ;
        RECT 102.525 157.955 103.275 158.475 ;
        RECT 100.205 157.185 100.535 157.815 ;
        RECT 100.705 157.015 100.915 157.835 ;
        RECT 103.445 157.785 104.195 158.305 ;
        RECT 101.605 157.015 101.895 157.740 ;
        RECT 102.525 157.015 104.195 157.785 ;
        RECT 104.365 157.690 104.535 158.490 ;
        RECT 104.820 158.465 105.485 158.635 ;
        RECT 105.835 158.635 106.005 159.395 ;
        RECT 106.185 158.805 106.515 159.565 ;
        RECT 105.835 158.465 106.500 158.635 ;
        RECT 106.685 158.490 106.955 159.395 ;
        RECT 104.820 158.320 104.990 158.465 ;
        RECT 104.705 157.990 104.990 158.320 ;
        RECT 106.330 158.320 106.500 158.465 ;
        RECT 104.820 157.735 104.990 157.990 ;
        RECT 105.225 157.915 105.555 158.285 ;
        RECT 105.765 157.915 106.095 158.285 ;
        RECT 106.330 157.990 106.615 158.320 ;
        RECT 106.330 157.735 106.500 157.990 ;
        RECT 104.365 157.185 104.625 157.690 ;
        RECT 104.820 157.565 105.485 157.735 ;
        RECT 104.805 157.015 105.135 157.395 ;
        RECT 105.315 157.185 105.485 157.565 ;
        RECT 105.835 157.565 106.500 157.735 ;
        RECT 106.785 157.690 106.955 158.490 ;
        RECT 105.835 157.185 106.005 157.565 ;
        RECT 106.185 157.015 106.515 157.395 ;
        RECT 106.695 157.185 106.955 157.690 ;
        RECT 108.045 158.425 108.385 159.395 ;
        RECT 108.555 158.425 108.725 159.565 ;
        RECT 108.995 158.765 109.245 159.565 ;
        RECT 109.890 158.595 110.220 159.395 ;
        RECT 110.520 158.765 110.850 159.565 ;
        RECT 111.020 158.595 111.350 159.395 ;
        RECT 108.915 158.425 111.350 158.595 ;
        RECT 112.645 158.475 116.155 159.565 ;
        RECT 116.440 158.935 116.725 159.395 ;
        RECT 116.895 159.105 117.165 159.565 ;
        RECT 116.440 158.715 117.395 158.935 ;
        RECT 108.045 157.815 108.220 158.425 ;
        RECT 108.915 158.175 109.085 158.425 ;
        RECT 108.390 158.005 109.085 158.175 ;
        RECT 109.260 158.005 109.680 158.205 ;
        RECT 109.850 158.005 110.180 158.205 ;
        RECT 110.350 158.005 110.680 158.205 ;
        RECT 108.045 157.185 108.385 157.815 ;
        RECT 108.555 157.015 108.805 157.815 ;
        RECT 108.995 157.665 110.220 157.835 ;
        RECT 108.995 157.185 109.325 157.665 ;
        RECT 109.495 157.015 109.720 157.475 ;
        RECT 109.890 157.185 110.220 157.665 ;
        RECT 110.850 157.795 111.020 158.425 ;
        RECT 111.205 158.005 111.555 158.255 ;
        RECT 112.645 157.955 114.335 158.475 ;
        RECT 110.850 157.185 111.350 157.795 ;
        RECT 114.505 157.785 116.155 158.305 ;
        RECT 116.325 157.985 117.015 158.545 ;
        RECT 117.185 157.815 117.395 158.715 ;
        RECT 112.645 157.015 116.155 157.785 ;
        RECT 116.440 157.645 117.395 157.815 ;
        RECT 117.565 158.545 117.965 159.395 ;
        RECT 118.155 158.935 118.435 159.395 ;
        RECT 118.955 159.105 119.280 159.565 ;
        RECT 118.155 158.715 119.280 158.935 ;
        RECT 117.565 157.985 118.660 158.545 ;
        RECT 118.830 158.255 119.280 158.715 ;
        RECT 119.450 158.425 119.835 159.395 ;
        RECT 120.930 159.130 126.275 159.565 ;
        RECT 116.440 157.185 116.725 157.645 ;
        RECT 116.895 157.015 117.165 157.475 ;
        RECT 117.565 157.185 117.965 157.985 ;
        RECT 118.830 157.925 119.385 158.255 ;
        RECT 118.830 157.815 119.280 157.925 ;
        RECT 118.155 157.645 119.280 157.815 ;
        RECT 119.555 157.755 119.835 158.425 ;
        RECT 122.520 157.880 122.870 159.130 ;
        RECT 126.445 158.475 127.655 159.565 ;
        RECT 118.155 157.185 118.435 157.645 ;
        RECT 118.955 157.015 119.280 157.475 ;
        RECT 119.450 157.185 119.835 157.755 ;
        RECT 124.350 157.560 124.690 158.390 ;
        RECT 126.445 157.935 126.965 158.475 ;
        RECT 127.135 157.765 127.655 158.305 ;
        RECT 120.930 157.015 126.275 157.560 ;
        RECT 126.445 157.015 127.655 157.765 ;
        RECT 14.580 156.845 127.740 157.015 ;
        RECT 14.665 156.095 15.875 156.845 ;
        RECT 17.340 156.505 17.595 156.665 ;
        RECT 17.255 156.335 17.595 156.505 ;
        RECT 17.775 156.385 18.060 156.845 ;
        RECT 17.340 156.135 17.595 156.335 ;
        RECT 14.665 155.555 15.185 156.095 ;
        RECT 15.355 155.385 15.875 155.925 ;
        RECT 14.665 154.295 15.875 155.385 ;
        RECT 17.340 155.275 17.520 156.135 ;
        RECT 18.240 155.935 18.490 156.585 ;
        RECT 17.690 155.605 18.490 155.935 ;
        RECT 17.340 154.605 17.595 155.275 ;
        RECT 17.775 154.295 18.060 155.095 ;
        RECT 18.240 155.015 18.490 155.605 ;
        RECT 18.690 156.250 19.010 156.580 ;
        RECT 19.190 156.365 19.850 156.845 ;
        RECT 20.050 156.455 20.900 156.625 ;
        RECT 18.690 155.355 18.880 156.250 ;
        RECT 19.200 155.925 19.860 156.195 ;
        RECT 19.530 155.865 19.860 155.925 ;
        RECT 19.050 155.695 19.380 155.755 ;
        RECT 20.050 155.695 20.220 156.455 ;
        RECT 21.460 156.385 21.780 156.845 ;
        RECT 21.980 156.205 22.230 156.635 ;
        RECT 22.520 156.405 22.930 156.845 ;
        RECT 23.100 156.465 24.115 156.665 ;
        RECT 20.390 156.035 21.640 156.205 ;
        RECT 20.390 155.915 20.720 156.035 ;
        RECT 19.050 155.525 20.950 155.695 ;
        RECT 18.690 155.185 20.610 155.355 ;
        RECT 18.690 155.165 19.010 155.185 ;
        RECT 18.240 154.505 18.570 155.015 ;
        RECT 18.840 154.555 19.010 155.165 ;
        RECT 20.780 155.015 20.950 155.525 ;
        RECT 21.120 155.455 21.300 155.865 ;
        RECT 21.470 155.275 21.640 156.035 ;
        RECT 19.180 154.295 19.510 154.985 ;
        RECT 19.740 154.845 20.950 155.015 ;
        RECT 21.120 154.965 21.640 155.275 ;
        RECT 21.810 155.865 22.230 156.205 ;
        RECT 22.520 155.865 22.930 156.195 ;
        RECT 21.810 155.095 22.000 155.865 ;
        RECT 23.100 155.735 23.270 156.465 ;
        RECT 24.415 156.295 24.585 156.625 ;
        RECT 24.755 156.465 25.085 156.845 ;
        RECT 23.440 155.915 23.790 156.285 ;
        RECT 23.100 155.695 23.520 155.735 ;
        RECT 22.170 155.525 23.520 155.695 ;
        RECT 22.170 155.365 22.420 155.525 ;
        RECT 22.930 155.095 23.180 155.355 ;
        RECT 21.810 154.845 23.180 155.095 ;
        RECT 19.740 154.555 19.980 154.845 ;
        RECT 20.780 154.765 20.950 154.845 ;
        RECT 20.180 154.295 20.600 154.675 ;
        RECT 20.780 154.515 21.410 154.765 ;
        RECT 21.880 154.295 22.210 154.675 ;
        RECT 22.380 154.555 22.550 154.845 ;
        RECT 23.350 154.680 23.520 155.525 ;
        RECT 23.970 155.355 24.190 156.225 ;
        RECT 24.415 156.105 25.110 156.295 ;
        RECT 23.690 154.975 24.190 155.355 ;
        RECT 24.360 155.305 24.770 155.925 ;
        RECT 24.940 155.135 25.110 156.105 ;
        RECT 24.415 154.965 25.110 155.135 ;
        RECT 22.730 154.295 23.110 154.675 ;
        RECT 23.350 154.510 24.180 154.680 ;
        RECT 24.415 154.465 24.585 154.965 ;
        RECT 24.755 154.295 25.085 154.795 ;
        RECT 25.300 154.465 25.525 156.585 ;
        RECT 25.695 156.465 26.025 156.845 ;
        RECT 26.195 156.295 26.365 156.585 ;
        RECT 25.700 156.125 26.365 156.295 ;
        RECT 26.625 156.170 26.885 156.675 ;
        RECT 27.065 156.465 27.395 156.845 ;
        RECT 27.575 156.295 27.745 156.675 ;
        RECT 25.700 155.135 25.930 156.125 ;
        RECT 26.100 155.305 26.450 155.955 ;
        RECT 26.625 155.370 26.795 156.170 ;
        RECT 27.080 156.125 27.745 156.295 ;
        RECT 27.080 155.870 27.250 156.125 ;
        RECT 28.005 156.095 29.215 156.845 ;
        RECT 26.965 155.540 27.250 155.870 ;
        RECT 27.485 155.575 27.815 155.945 ;
        RECT 27.080 155.395 27.250 155.540 ;
        RECT 25.700 154.965 26.365 155.135 ;
        RECT 25.695 154.295 26.025 154.795 ;
        RECT 26.195 154.465 26.365 154.965 ;
        RECT 26.625 154.465 26.895 155.370 ;
        RECT 27.080 155.225 27.745 155.395 ;
        RECT 27.065 154.295 27.395 155.055 ;
        RECT 27.575 154.465 27.745 155.225 ;
        RECT 28.005 155.385 28.525 155.925 ;
        RECT 28.695 155.555 29.215 156.095 ;
        RECT 29.385 156.075 32.895 156.845 ;
        RECT 29.385 155.385 31.075 155.905 ;
        RECT 31.245 155.555 32.895 156.075 ;
        RECT 33.340 156.035 33.585 156.640 ;
        RECT 33.805 156.310 34.315 156.845 ;
        RECT 33.065 155.865 34.295 156.035 ;
        RECT 28.005 154.295 29.215 155.385 ;
        RECT 29.385 154.295 32.895 155.385 ;
        RECT 33.065 155.055 33.405 155.865 ;
        RECT 33.575 155.300 34.325 155.490 ;
        RECT 33.065 154.645 33.580 155.055 ;
        RECT 33.815 154.295 33.985 155.055 ;
        RECT 34.155 154.635 34.325 155.300 ;
        RECT 34.495 155.315 34.685 156.675 ;
        RECT 34.855 156.505 35.130 156.675 ;
        RECT 34.855 156.335 35.135 156.505 ;
        RECT 34.855 155.515 35.130 156.335 ;
        RECT 35.320 156.310 35.850 156.675 ;
        RECT 36.275 156.445 36.605 156.845 ;
        RECT 35.675 156.275 35.850 156.310 ;
        RECT 35.335 155.315 35.505 156.115 ;
        RECT 34.495 155.145 35.505 155.315 ;
        RECT 35.675 156.105 36.605 156.275 ;
        RECT 36.775 156.105 37.030 156.675 ;
        RECT 37.205 156.120 37.495 156.845 ;
        RECT 35.675 154.975 35.845 156.105 ;
        RECT 36.435 155.935 36.605 156.105 ;
        RECT 34.720 154.805 35.845 154.975 ;
        RECT 36.015 155.605 36.210 155.935 ;
        RECT 36.435 155.605 36.690 155.935 ;
        RECT 36.015 154.635 36.185 155.605 ;
        RECT 36.860 155.435 37.030 156.105 ;
        RECT 38.125 156.075 39.795 156.845 ;
        RECT 34.155 154.465 36.185 154.635 ;
        RECT 36.355 154.295 36.525 155.435 ;
        RECT 36.695 154.465 37.030 155.435 ;
        RECT 37.205 154.295 37.495 155.460 ;
        RECT 38.125 155.385 38.875 155.905 ;
        RECT 39.045 155.555 39.795 156.075 ;
        RECT 39.965 156.045 40.305 156.675 ;
        RECT 40.475 156.045 40.725 156.845 ;
        RECT 40.915 156.195 41.245 156.675 ;
        RECT 41.415 156.385 41.640 156.845 ;
        RECT 41.810 156.195 42.140 156.675 ;
        RECT 39.965 155.435 40.140 156.045 ;
        RECT 40.915 156.025 42.140 156.195 ;
        RECT 42.770 156.065 43.270 156.675 ;
        RECT 40.310 155.685 41.005 155.855 ;
        RECT 40.835 155.435 41.005 155.685 ;
        RECT 41.180 155.655 41.600 155.855 ;
        RECT 41.770 155.655 42.100 155.855 ;
        RECT 42.270 155.655 42.600 155.855 ;
        RECT 42.770 155.435 42.940 156.065 ;
        RECT 43.645 156.045 43.985 156.675 ;
        RECT 44.155 156.045 44.405 156.845 ;
        RECT 44.595 156.195 44.925 156.675 ;
        RECT 45.095 156.385 45.320 156.845 ;
        RECT 45.490 156.195 45.820 156.675 ;
        RECT 43.125 155.605 43.475 155.855 ;
        RECT 43.645 155.435 43.820 156.045 ;
        RECT 44.595 156.025 45.820 156.195 ;
        RECT 46.450 156.065 46.950 156.675 ;
        RECT 43.990 155.685 44.685 155.855 ;
        RECT 44.515 155.435 44.685 155.685 ;
        RECT 44.860 155.655 45.280 155.855 ;
        RECT 45.450 155.655 45.780 155.855 ;
        RECT 45.950 155.655 46.280 155.855 ;
        RECT 46.450 155.435 46.620 156.065 ;
        RECT 47.325 156.045 47.665 156.675 ;
        RECT 47.835 156.045 48.085 156.845 ;
        RECT 48.275 156.195 48.605 156.675 ;
        RECT 48.775 156.385 49.000 156.845 ;
        RECT 49.170 156.195 49.500 156.675 ;
        RECT 46.805 155.605 47.155 155.855 ;
        RECT 47.325 155.435 47.500 156.045 ;
        RECT 48.275 156.025 49.500 156.195 ;
        RECT 50.130 156.065 50.630 156.675 ;
        RECT 51.465 156.075 53.135 156.845 ;
        RECT 47.670 155.685 48.365 155.855 ;
        RECT 48.195 155.435 48.365 155.685 ;
        RECT 48.540 155.655 48.960 155.855 ;
        RECT 49.130 155.655 49.460 155.855 ;
        RECT 49.630 155.655 49.960 155.855 ;
        RECT 50.130 155.435 50.300 156.065 ;
        RECT 50.485 155.605 50.835 155.855 ;
        RECT 38.125 154.295 39.795 155.385 ;
        RECT 39.965 154.465 40.305 155.435 ;
        RECT 40.475 154.295 40.645 155.435 ;
        RECT 40.835 155.265 43.270 155.435 ;
        RECT 40.915 154.295 41.165 155.095 ;
        RECT 41.810 154.465 42.140 155.265 ;
        RECT 42.440 154.295 42.770 155.095 ;
        RECT 42.940 154.465 43.270 155.265 ;
        RECT 43.645 154.465 43.985 155.435 ;
        RECT 44.155 154.295 44.325 155.435 ;
        RECT 44.515 155.265 46.950 155.435 ;
        RECT 44.595 154.295 44.845 155.095 ;
        RECT 45.490 154.465 45.820 155.265 ;
        RECT 46.120 154.295 46.450 155.095 ;
        RECT 46.620 154.465 46.950 155.265 ;
        RECT 47.325 154.465 47.665 155.435 ;
        RECT 47.835 154.295 48.005 155.435 ;
        RECT 48.195 155.265 50.630 155.435 ;
        RECT 48.275 154.295 48.525 155.095 ;
        RECT 49.170 154.465 49.500 155.265 ;
        RECT 49.800 154.295 50.130 155.095 ;
        RECT 50.300 154.465 50.630 155.265 ;
        RECT 51.465 155.385 52.215 155.905 ;
        RECT 52.385 155.555 53.135 156.075 ;
        RECT 53.680 156.135 53.935 156.665 ;
        RECT 54.115 156.385 54.400 156.845 ;
        RECT 51.465 154.295 53.135 155.385 ;
        RECT 53.680 155.275 53.860 156.135 ;
        RECT 54.580 155.935 54.830 156.585 ;
        RECT 54.030 155.605 54.830 155.935 ;
        RECT 53.680 154.805 53.935 155.275 ;
        RECT 53.595 154.635 53.935 154.805 ;
        RECT 53.680 154.605 53.935 154.635 ;
        RECT 54.115 154.295 54.400 155.095 ;
        RECT 54.580 155.015 54.830 155.605 ;
        RECT 55.030 156.250 55.350 156.580 ;
        RECT 55.530 156.365 56.190 156.845 ;
        RECT 56.390 156.455 57.240 156.625 ;
        RECT 55.030 155.355 55.220 156.250 ;
        RECT 55.540 155.925 56.200 156.195 ;
        RECT 55.870 155.865 56.200 155.925 ;
        RECT 55.390 155.695 55.720 155.755 ;
        RECT 56.390 155.695 56.560 156.455 ;
        RECT 57.800 156.385 58.120 156.845 ;
        RECT 58.320 156.205 58.570 156.635 ;
        RECT 58.860 156.405 59.270 156.845 ;
        RECT 59.440 156.465 60.455 156.665 ;
        RECT 56.730 156.035 57.980 156.205 ;
        RECT 56.730 155.915 57.060 156.035 ;
        RECT 55.390 155.525 57.290 155.695 ;
        RECT 55.030 155.185 56.950 155.355 ;
        RECT 55.030 155.165 55.350 155.185 ;
        RECT 54.580 154.505 54.910 155.015 ;
        RECT 55.180 154.555 55.350 155.165 ;
        RECT 57.120 155.015 57.290 155.525 ;
        RECT 57.460 155.455 57.640 155.865 ;
        RECT 57.810 155.275 57.980 156.035 ;
        RECT 55.520 154.295 55.850 154.985 ;
        RECT 56.080 154.845 57.290 155.015 ;
        RECT 57.460 154.965 57.980 155.275 ;
        RECT 58.150 155.865 58.570 156.205 ;
        RECT 58.860 155.865 59.270 156.195 ;
        RECT 58.150 155.095 58.340 155.865 ;
        RECT 59.440 155.735 59.610 156.465 ;
        RECT 60.755 156.295 60.925 156.625 ;
        RECT 61.095 156.465 61.425 156.845 ;
        RECT 59.780 155.915 60.130 156.285 ;
        RECT 59.440 155.695 59.860 155.735 ;
        RECT 58.510 155.525 59.860 155.695 ;
        RECT 58.510 155.365 58.760 155.525 ;
        RECT 59.270 155.095 59.520 155.355 ;
        RECT 58.150 154.845 59.520 155.095 ;
        RECT 56.080 154.555 56.320 154.845 ;
        RECT 57.120 154.765 57.290 154.845 ;
        RECT 56.520 154.295 56.940 154.675 ;
        RECT 57.120 154.515 57.750 154.765 ;
        RECT 58.220 154.295 58.550 154.675 ;
        RECT 58.720 154.555 58.890 154.845 ;
        RECT 59.690 154.680 59.860 155.525 ;
        RECT 60.310 155.355 60.530 156.225 ;
        RECT 60.755 156.105 61.450 156.295 ;
        RECT 60.030 154.975 60.530 155.355 ;
        RECT 60.700 155.305 61.110 155.925 ;
        RECT 61.280 155.135 61.450 156.105 ;
        RECT 60.755 154.965 61.450 155.135 ;
        RECT 59.070 154.295 59.450 154.675 ;
        RECT 59.690 154.510 60.520 154.680 ;
        RECT 60.755 154.465 60.925 154.965 ;
        RECT 61.095 154.295 61.425 154.795 ;
        RECT 61.640 154.465 61.865 156.585 ;
        RECT 62.035 156.465 62.365 156.845 ;
        RECT 62.535 156.295 62.705 156.585 ;
        RECT 62.040 156.125 62.705 156.295 ;
        RECT 62.040 155.135 62.270 156.125 ;
        RECT 62.965 156.120 63.255 156.845 ;
        RECT 63.885 156.075 65.555 156.845 ;
        RECT 65.815 156.365 66.115 156.845 ;
        RECT 66.285 156.195 66.545 156.650 ;
        RECT 66.715 156.365 66.975 156.845 ;
        RECT 67.155 156.195 67.415 156.650 ;
        RECT 67.585 156.365 67.835 156.845 ;
        RECT 68.015 156.195 68.275 156.650 ;
        RECT 68.445 156.365 68.695 156.845 ;
        RECT 68.875 156.195 69.135 156.650 ;
        RECT 69.305 156.365 69.550 156.845 ;
        RECT 69.720 156.195 69.995 156.650 ;
        RECT 70.165 156.365 70.410 156.845 ;
        RECT 70.580 156.195 70.840 156.650 ;
        RECT 71.010 156.365 71.270 156.845 ;
        RECT 71.440 156.195 71.700 156.650 ;
        RECT 71.870 156.365 72.130 156.845 ;
        RECT 72.300 156.195 72.560 156.650 ;
        RECT 72.730 156.285 72.990 156.845 ;
        RECT 62.440 155.305 62.790 155.955 ;
        RECT 62.040 154.965 62.705 155.135 ;
        RECT 62.035 154.295 62.365 154.795 ;
        RECT 62.535 154.465 62.705 154.965 ;
        RECT 62.965 154.295 63.255 155.460 ;
        RECT 63.885 155.385 64.635 155.905 ;
        RECT 64.805 155.555 65.555 156.075 ;
        RECT 65.815 156.025 72.560 156.195 ;
        RECT 65.815 155.485 66.980 156.025 ;
        RECT 73.160 155.855 73.410 156.665 ;
        RECT 73.590 156.320 73.850 156.845 ;
        RECT 74.020 155.855 74.270 156.665 ;
        RECT 74.450 156.335 74.755 156.845 ;
        RECT 67.150 155.605 74.270 155.855 ;
        RECT 74.440 155.605 74.755 156.165 ;
        RECT 74.925 156.075 76.595 156.845 ;
        RECT 65.785 155.435 66.980 155.485 ;
        RECT 63.885 154.295 65.555 155.385 ;
        RECT 65.785 155.315 72.560 155.435 ;
        RECT 65.815 155.210 72.560 155.315 ;
        RECT 65.815 154.295 66.085 155.040 ;
        RECT 66.255 154.470 66.545 155.210 ;
        RECT 67.155 155.195 72.560 155.210 ;
        RECT 66.715 154.300 66.970 155.025 ;
        RECT 67.155 154.470 67.415 155.195 ;
        RECT 67.585 154.300 67.830 155.025 ;
        RECT 68.015 154.470 68.275 155.195 ;
        RECT 68.445 154.300 68.690 155.025 ;
        RECT 68.875 154.470 69.135 155.195 ;
        RECT 69.305 154.300 69.550 155.025 ;
        RECT 69.720 154.470 69.980 155.195 ;
        RECT 70.150 154.300 70.410 155.025 ;
        RECT 70.580 154.470 70.840 155.195 ;
        RECT 71.010 154.300 71.270 155.025 ;
        RECT 71.440 154.470 71.700 155.195 ;
        RECT 71.870 154.300 72.130 155.025 ;
        RECT 72.300 154.470 72.560 155.195 ;
        RECT 72.730 154.300 72.990 155.095 ;
        RECT 73.160 154.470 73.410 155.605 ;
        RECT 66.715 154.295 72.990 154.300 ;
        RECT 73.590 154.295 73.850 155.105 ;
        RECT 74.025 154.465 74.270 155.605 ;
        RECT 74.925 155.385 75.675 155.905 ;
        RECT 75.845 155.555 76.595 156.075 ;
        RECT 76.765 156.045 77.105 156.675 ;
        RECT 77.275 156.045 77.525 156.845 ;
        RECT 77.715 156.195 78.045 156.675 ;
        RECT 78.215 156.385 78.440 156.845 ;
        RECT 78.610 156.195 78.940 156.675 ;
        RECT 76.765 155.435 76.940 156.045 ;
        RECT 77.715 156.025 78.940 156.195 ;
        RECT 79.570 156.065 80.070 156.675 ;
        RECT 77.110 155.685 77.805 155.855 ;
        RECT 77.635 155.435 77.805 155.685 ;
        RECT 77.980 155.655 78.400 155.855 ;
        RECT 78.570 155.655 78.900 155.855 ;
        RECT 79.070 155.655 79.400 155.855 ;
        RECT 79.570 155.435 79.740 156.065 ;
        RECT 80.445 156.045 80.785 156.675 ;
        RECT 80.955 156.045 81.205 156.845 ;
        RECT 81.395 156.195 81.725 156.675 ;
        RECT 81.895 156.385 82.120 156.845 ;
        RECT 82.290 156.195 82.620 156.675 ;
        RECT 79.925 155.605 80.275 155.855 ;
        RECT 80.445 155.435 80.620 156.045 ;
        RECT 81.395 156.025 82.620 156.195 ;
        RECT 83.250 156.065 83.750 156.675 ;
        RECT 85.045 156.075 88.555 156.845 ;
        RECT 88.725 156.120 89.015 156.845 ;
        RECT 89.185 156.075 91.775 156.845 ;
        RECT 91.950 156.300 97.295 156.845 ;
        RECT 80.790 155.685 81.485 155.855 ;
        RECT 81.315 155.435 81.485 155.685 ;
        RECT 81.660 155.655 82.080 155.855 ;
        RECT 82.250 155.655 82.580 155.855 ;
        RECT 82.750 155.655 83.080 155.855 ;
        RECT 83.250 155.435 83.420 156.065 ;
        RECT 83.605 155.605 83.955 155.855 ;
        RECT 74.450 154.295 74.745 155.105 ;
        RECT 74.925 154.295 76.595 155.385 ;
        RECT 76.765 154.465 77.105 155.435 ;
        RECT 77.275 154.295 77.445 155.435 ;
        RECT 77.635 155.265 80.070 155.435 ;
        RECT 77.715 154.295 77.965 155.095 ;
        RECT 78.610 154.465 78.940 155.265 ;
        RECT 79.240 154.295 79.570 155.095 ;
        RECT 79.740 154.465 80.070 155.265 ;
        RECT 80.445 154.465 80.785 155.435 ;
        RECT 80.955 154.295 81.125 155.435 ;
        RECT 81.315 155.265 83.750 155.435 ;
        RECT 81.395 154.295 81.645 155.095 ;
        RECT 82.290 154.465 82.620 155.265 ;
        RECT 82.920 154.295 83.250 155.095 ;
        RECT 83.420 154.465 83.750 155.265 ;
        RECT 85.045 155.385 86.735 155.905 ;
        RECT 86.905 155.555 88.555 156.075 ;
        RECT 85.045 154.295 88.555 155.385 ;
        RECT 88.725 154.295 89.015 155.460 ;
        RECT 89.185 155.385 90.395 155.905 ;
        RECT 90.565 155.555 91.775 156.075 ;
        RECT 89.185 154.295 91.775 155.385 ;
        RECT 93.540 154.730 93.890 155.980 ;
        RECT 95.370 155.470 95.710 156.300 ;
        RECT 97.670 156.065 98.170 156.675 ;
        RECT 97.465 155.605 97.815 155.855 ;
        RECT 98.000 155.435 98.170 156.065 ;
        RECT 98.800 156.195 99.130 156.675 ;
        RECT 99.300 156.385 99.525 156.845 ;
        RECT 99.695 156.195 100.025 156.675 ;
        RECT 98.800 156.025 100.025 156.195 ;
        RECT 100.215 156.045 100.465 156.845 ;
        RECT 100.635 156.045 100.975 156.675 ;
        RECT 101.605 156.075 103.275 156.845 ;
        RECT 98.340 155.655 98.670 155.855 ;
        RECT 98.840 155.655 99.170 155.855 ;
        RECT 99.340 155.655 99.760 155.855 ;
        RECT 99.935 155.685 100.630 155.855 ;
        RECT 99.935 155.435 100.105 155.685 ;
        RECT 100.800 155.435 100.975 156.045 ;
        RECT 97.670 155.265 100.105 155.435 ;
        RECT 91.950 154.295 97.295 154.730 ;
        RECT 97.670 154.465 98.000 155.265 ;
        RECT 98.170 154.295 98.500 155.095 ;
        RECT 98.800 154.465 99.130 155.265 ;
        RECT 99.775 154.295 100.025 155.095 ;
        RECT 100.295 154.295 100.465 155.435 ;
        RECT 100.635 154.465 100.975 155.435 ;
        RECT 101.605 155.385 102.355 155.905 ;
        RECT 102.525 155.555 103.275 156.075 ;
        RECT 103.445 156.045 103.785 156.675 ;
        RECT 103.955 156.045 104.205 156.845 ;
        RECT 104.395 156.195 104.725 156.675 ;
        RECT 104.895 156.385 105.120 156.845 ;
        RECT 105.290 156.195 105.620 156.675 ;
        RECT 103.445 155.435 103.620 156.045 ;
        RECT 104.395 156.025 105.620 156.195 ;
        RECT 106.250 156.065 106.750 156.675 ;
        RECT 107.330 156.065 107.830 156.675 ;
        RECT 103.790 155.685 104.485 155.855 ;
        RECT 104.315 155.435 104.485 155.685 ;
        RECT 104.660 155.655 105.080 155.855 ;
        RECT 105.250 155.655 105.580 155.855 ;
        RECT 105.750 155.655 106.080 155.855 ;
        RECT 106.250 155.435 106.420 156.065 ;
        RECT 106.605 155.605 106.955 155.855 ;
        RECT 107.125 155.605 107.475 155.855 ;
        RECT 107.660 155.435 107.830 156.065 ;
        RECT 108.460 156.195 108.790 156.675 ;
        RECT 108.960 156.385 109.185 156.845 ;
        RECT 109.355 156.195 109.685 156.675 ;
        RECT 108.460 156.025 109.685 156.195 ;
        RECT 109.875 156.045 110.125 156.845 ;
        RECT 110.295 156.045 110.635 156.675 ;
        RECT 110.805 156.075 114.315 156.845 ;
        RECT 114.485 156.120 114.775 156.845 ;
        RECT 114.945 156.095 116.155 156.845 ;
        RECT 108.000 155.655 108.330 155.855 ;
        RECT 108.500 155.655 108.830 155.855 ;
        RECT 109.000 155.655 109.420 155.855 ;
        RECT 109.595 155.685 110.290 155.855 ;
        RECT 109.595 155.435 109.765 155.685 ;
        RECT 110.460 155.435 110.635 156.045 ;
        RECT 101.605 154.295 103.275 155.385 ;
        RECT 103.445 154.465 103.785 155.435 ;
        RECT 103.955 154.295 104.125 155.435 ;
        RECT 104.315 155.265 106.750 155.435 ;
        RECT 104.395 154.295 104.645 155.095 ;
        RECT 105.290 154.465 105.620 155.265 ;
        RECT 105.920 154.295 106.250 155.095 ;
        RECT 106.420 154.465 106.750 155.265 ;
        RECT 107.330 155.265 109.765 155.435 ;
        RECT 107.330 154.465 107.660 155.265 ;
        RECT 107.830 154.295 108.160 155.095 ;
        RECT 108.460 154.465 108.790 155.265 ;
        RECT 109.435 154.295 109.685 155.095 ;
        RECT 109.955 154.295 110.125 155.435 ;
        RECT 110.295 154.465 110.635 155.435 ;
        RECT 110.805 155.385 112.495 155.905 ;
        RECT 112.665 155.555 114.315 156.075 ;
        RECT 110.805 154.295 114.315 155.385 ;
        RECT 114.485 154.295 114.775 155.460 ;
        RECT 114.945 155.385 115.465 155.925 ;
        RECT 115.635 155.555 116.155 156.095 ;
        RECT 116.415 156.195 116.585 156.675 ;
        RECT 116.765 156.365 117.005 156.845 ;
        RECT 117.255 156.195 117.425 156.675 ;
        RECT 117.595 156.365 117.925 156.845 ;
        RECT 118.095 156.195 118.265 156.675 ;
        RECT 116.415 156.025 117.050 156.195 ;
        RECT 117.255 156.025 118.265 156.195 ;
        RECT 118.435 156.045 118.765 156.845 ;
        RECT 119.085 156.075 120.755 156.845 ;
        RECT 120.930 156.300 126.275 156.845 ;
        RECT 116.880 155.855 117.050 156.025 ;
        RECT 116.330 155.615 116.710 155.855 ;
        RECT 116.880 155.685 117.380 155.855 ;
        RECT 116.880 155.445 117.050 155.685 ;
        RECT 117.770 155.485 118.265 156.025 ;
        RECT 114.945 154.295 116.155 155.385 ;
        RECT 116.335 155.275 117.050 155.445 ;
        RECT 117.255 155.315 118.265 155.485 ;
        RECT 116.335 154.465 116.665 155.275 ;
        RECT 116.835 154.295 117.075 155.095 ;
        RECT 117.255 154.465 117.425 155.315 ;
        RECT 117.595 154.295 117.925 155.095 ;
        RECT 118.095 154.465 118.265 155.315 ;
        RECT 118.435 154.295 118.765 155.445 ;
        RECT 119.085 155.385 119.835 155.905 ;
        RECT 120.005 155.555 120.755 156.075 ;
        RECT 119.085 154.295 120.755 155.385 ;
        RECT 122.520 154.730 122.870 155.980 ;
        RECT 124.350 155.470 124.690 156.300 ;
        RECT 126.445 156.095 127.655 156.845 ;
        RECT 126.445 155.385 126.965 155.925 ;
        RECT 127.135 155.555 127.655 156.095 ;
        RECT 120.930 154.295 126.275 154.730 ;
        RECT 126.445 154.295 127.655 155.385 ;
        RECT 14.580 154.125 127.740 154.295 ;
        RECT 14.665 153.035 15.875 154.125 ;
        RECT 14.665 152.325 15.185 152.865 ;
        RECT 15.355 152.495 15.875 153.035 ;
        RECT 16.505 153.035 20.015 154.125 ;
        RECT 20.185 153.365 20.700 153.775 ;
        RECT 20.935 153.365 21.105 154.125 ;
        RECT 21.275 153.785 23.305 153.955 ;
        RECT 16.505 152.515 18.195 153.035 ;
        RECT 18.365 152.345 20.015 152.865 ;
        RECT 20.185 152.555 20.525 153.365 ;
        RECT 21.275 153.120 21.445 153.785 ;
        RECT 21.840 153.445 22.965 153.615 ;
        RECT 20.695 152.930 21.445 153.120 ;
        RECT 21.615 153.105 22.625 153.275 ;
        RECT 20.185 152.385 21.415 152.555 ;
        RECT 14.665 151.575 15.875 152.325 ;
        RECT 16.505 151.575 20.015 152.345 ;
        RECT 20.460 151.780 20.705 152.385 ;
        RECT 20.925 151.575 21.435 152.110 ;
        RECT 21.615 151.745 21.805 153.105 ;
        RECT 21.975 152.085 22.250 152.905 ;
        RECT 22.455 152.305 22.625 153.105 ;
        RECT 22.795 152.315 22.965 153.445 ;
        RECT 23.135 152.815 23.305 153.785 ;
        RECT 23.475 152.985 23.645 154.125 ;
        RECT 23.815 152.985 24.150 153.955 ;
        RECT 23.135 152.485 23.330 152.815 ;
        RECT 23.555 152.485 23.810 152.815 ;
        RECT 23.555 152.315 23.725 152.485 ;
        RECT 23.980 152.315 24.150 152.985 ;
        RECT 24.325 152.960 24.615 154.125 ;
        RECT 24.785 153.035 25.995 154.125 ;
        RECT 26.165 153.035 29.675 154.125 ;
        RECT 30.220 153.145 30.475 153.815 ;
        RECT 30.655 153.325 30.940 154.125 ;
        RECT 31.120 153.405 31.450 153.915 ;
        RECT 24.785 152.495 25.305 153.035 ;
        RECT 25.475 152.325 25.995 152.865 ;
        RECT 26.165 152.515 27.855 153.035 ;
        RECT 28.025 152.345 29.675 152.865 ;
        RECT 22.795 152.145 23.725 152.315 ;
        RECT 22.795 152.110 22.970 152.145 ;
        RECT 21.975 151.915 22.255 152.085 ;
        RECT 21.975 151.745 22.250 151.915 ;
        RECT 22.440 151.745 22.970 152.110 ;
        RECT 23.395 151.575 23.725 151.975 ;
        RECT 23.895 151.745 24.150 152.315 ;
        RECT 24.325 151.575 24.615 152.300 ;
        RECT 24.785 151.575 25.995 152.325 ;
        RECT 26.165 151.575 29.675 152.345 ;
        RECT 30.220 152.285 30.400 153.145 ;
        RECT 31.120 152.815 31.370 153.405 ;
        RECT 31.720 153.255 31.890 153.865 ;
        RECT 32.060 153.435 32.390 154.125 ;
        RECT 32.620 153.575 32.860 153.865 ;
        RECT 33.060 153.745 33.480 154.125 ;
        RECT 33.660 153.655 34.290 153.905 ;
        RECT 34.760 153.745 35.090 154.125 ;
        RECT 33.660 153.575 33.830 153.655 ;
        RECT 35.260 153.575 35.430 153.865 ;
        RECT 35.610 153.745 35.990 154.125 ;
        RECT 36.230 153.740 37.060 153.910 ;
        RECT 32.620 153.405 33.830 153.575 ;
        RECT 30.570 152.485 31.370 152.815 ;
        RECT 30.220 152.085 30.475 152.285 ;
        RECT 30.135 151.915 30.475 152.085 ;
        RECT 30.220 151.755 30.475 151.915 ;
        RECT 30.655 151.575 30.940 152.035 ;
        RECT 31.120 151.835 31.370 152.485 ;
        RECT 31.570 153.235 31.890 153.255 ;
        RECT 31.570 153.065 33.490 153.235 ;
        RECT 31.570 152.170 31.760 153.065 ;
        RECT 33.660 152.895 33.830 153.405 ;
        RECT 34.000 153.145 34.520 153.455 ;
        RECT 31.930 152.725 33.830 152.895 ;
        RECT 31.930 152.665 32.260 152.725 ;
        RECT 32.410 152.495 32.740 152.555 ;
        RECT 32.080 152.225 32.740 152.495 ;
        RECT 31.570 151.840 31.890 152.170 ;
        RECT 32.070 151.575 32.730 152.055 ;
        RECT 32.930 151.965 33.100 152.725 ;
        RECT 34.000 152.555 34.180 152.965 ;
        RECT 33.270 152.385 33.600 152.505 ;
        RECT 34.350 152.385 34.520 153.145 ;
        RECT 33.270 152.215 34.520 152.385 ;
        RECT 34.690 153.325 36.060 153.575 ;
        RECT 34.690 152.555 34.880 153.325 ;
        RECT 35.810 153.065 36.060 153.325 ;
        RECT 35.050 152.895 35.300 153.055 ;
        RECT 36.230 152.895 36.400 153.740 ;
        RECT 37.295 153.455 37.465 153.955 ;
        RECT 37.635 153.625 37.965 154.125 ;
        RECT 36.570 153.065 37.070 153.445 ;
        RECT 37.295 153.285 37.990 153.455 ;
        RECT 35.050 152.725 36.400 152.895 ;
        RECT 35.980 152.685 36.400 152.725 ;
        RECT 34.690 152.215 35.110 152.555 ;
        RECT 35.400 152.225 35.810 152.555 ;
        RECT 32.930 151.795 33.780 151.965 ;
        RECT 34.340 151.575 34.660 152.035 ;
        RECT 34.860 151.785 35.110 152.215 ;
        RECT 35.400 151.575 35.810 152.015 ;
        RECT 35.980 151.955 36.150 152.685 ;
        RECT 36.320 152.135 36.670 152.505 ;
        RECT 36.850 152.195 37.070 153.065 ;
        RECT 37.240 152.495 37.650 153.115 ;
        RECT 37.820 152.315 37.990 153.285 ;
        RECT 37.295 152.125 37.990 152.315 ;
        RECT 35.980 151.755 36.995 151.955 ;
        RECT 37.295 151.795 37.465 152.125 ;
        RECT 37.635 151.575 37.965 151.955 ;
        RECT 38.180 151.835 38.405 153.955 ;
        RECT 38.575 153.625 38.905 154.125 ;
        RECT 39.075 153.455 39.245 153.955 ;
        RECT 38.580 153.285 39.245 153.455 ;
        RECT 38.580 152.295 38.810 153.285 ;
        RECT 38.980 152.465 39.330 153.115 ;
        RECT 39.505 152.985 39.845 153.955 ;
        RECT 40.015 152.985 40.185 154.125 ;
        RECT 40.455 153.325 40.705 154.125 ;
        RECT 41.350 153.155 41.680 153.955 ;
        RECT 41.980 153.325 42.310 154.125 ;
        RECT 42.480 153.155 42.810 153.955 ;
        RECT 40.375 152.985 42.810 153.155 ;
        RECT 43.185 153.035 44.395 154.125 ;
        RECT 44.570 153.690 49.915 154.125 ;
        RECT 39.505 152.375 39.680 152.985 ;
        RECT 40.375 152.735 40.545 152.985 ;
        RECT 39.850 152.565 40.545 152.735 ;
        RECT 40.720 152.565 41.140 152.765 ;
        RECT 41.310 152.565 41.640 152.765 ;
        RECT 41.810 152.565 42.140 152.765 ;
        RECT 38.580 152.125 39.245 152.295 ;
        RECT 38.575 151.575 38.905 151.955 ;
        RECT 39.075 151.835 39.245 152.125 ;
        RECT 39.505 151.745 39.845 152.375 ;
        RECT 40.015 151.575 40.265 152.375 ;
        RECT 40.455 152.225 41.680 152.395 ;
        RECT 40.455 151.745 40.785 152.225 ;
        RECT 40.955 151.575 41.180 152.035 ;
        RECT 41.350 151.745 41.680 152.225 ;
        RECT 42.310 152.355 42.480 152.985 ;
        RECT 42.665 152.565 43.015 152.815 ;
        RECT 43.185 152.495 43.705 153.035 ;
        RECT 42.310 151.745 42.810 152.355 ;
        RECT 43.875 152.325 44.395 152.865 ;
        RECT 46.160 152.440 46.510 153.690 ;
        RECT 50.085 152.960 50.375 154.125 ;
        RECT 51.470 153.690 56.815 154.125 ;
        RECT 43.185 151.575 44.395 152.325 ;
        RECT 47.990 152.120 48.330 152.950 ;
        RECT 53.060 152.440 53.410 153.690 ;
        RECT 57.025 152.985 57.255 154.125 ;
        RECT 57.425 152.975 57.755 153.955 ;
        RECT 57.925 152.985 58.135 154.125 ;
        RECT 58.740 153.145 58.995 153.815 ;
        RECT 59.175 153.325 59.460 154.125 ;
        RECT 59.640 153.405 59.970 153.915 ;
        RECT 44.570 151.575 49.915 152.120 ;
        RECT 50.085 151.575 50.375 152.300 ;
        RECT 54.890 152.120 55.230 152.950 ;
        RECT 57.005 152.565 57.335 152.815 ;
        RECT 51.470 151.575 56.815 152.120 ;
        RECT 57.025 151.575 57.255 152.395 ;
        RECT 57.505 152.375 57.755 152.975 ;
        RECT 57.425 151.745 57.755 152.375 ;
        RECT 57.925 151.575 58.135 152.395 ;
        RECT 58.740 152.285 58.920 153.145 ;
        RECT 59.640 152.815 59.890 153.405 ;
        RECT 60.240 153.255 60.410 153.865 ;
        RECT 60.580 153.435 60.910 154.125 ;
        RECT 61.140 153.575 61.380 153.865 ;
        RECT 61.580 153.745 62.000 154.125 ;
        RECT 62.180 153.655 62.810 153.905 ;
        RECT 63.280 153.745 63.610 154.125 ;
        RECT 62.180 153.575 62.350 153.655 ;
        RECT 63.780 153.575 63.950 153.865 ;
        RECT 64.130 153.745 64.510 154.125 ;
        RECT 64.750 153.740 65.580 153.910 ;
        RECT 61.140 153.405 62.350 153.575 ;
        RECT 59.090 152.485 59.890 152.815 ;
        RECT 58.740 152.085 58.995 152.285 ;
        RECT 58.655 151.915 58.995 152.085 ;
        RECT 58.740 151.755 58.995 151.915 ;
        RECT 59.175 151.575 59.460 152.035 ;
        RECT 59.640 151.835 59.890 152.485 ;
        RECT 60.090 153.235 60.410 153.255 ;
        RECT 60.090 153.065 62.010 153.235 ;
        RECT 60.090 152.170 60.280 153.065 ;
        RECT 62.180 152.895 62.350 153.405 ;
        RECT 62.520 153.145 63.040 153.455 ;
        RECT 60.450 152.725 62.350 152.895 ;
        RECT 60.450 152.665 60.780 152.725 ;
        RECT 60.930 152.495 61.260 152.555 ;
        RECT 60.600 152.225 61.260 152.495 ;
        RECT 60.090 151.840 60.410 152.170 ;
        RECT 60.590 151.575 61.250 152.055 ;
        RECT 61.450 151.965 61.620 152.725 ;
        RECT 62.520 152.555 62.700 152.965 ;
        RECT 61.790 152.385 62.120 152.505 ;
        RECT 62.870 152.385 63.040 153.145 ;
        RECT 61.790 152.215 63.040 152.385 ;
        RECT 63.210 153.325 64.580 153.575 ;
        RECT 63.210 152.555 63.400 153.325 ;
        RECT 64.330 153.065 64.580 153.325 ;
        RECT 63.570 152.895 63.820 153.055 ;
        RECT 64.750 152.895 64.920 153.740 ;
        RECT 65.815 153.455 65.985 153.955 ;
        RECT 66.155 153.625 66.485 154.125 ;
        RECT 65.090 153.065 65.590 153.445 ;
        RECT 65.815 153.285 66.510 153.455 ;
        RECT 63.570 152.725 64.920 152.895 ;
        RECT 64.500 152.685 64.920 152.725 ;
        RECT 63.210 152.215 63.630 152.555 ;
        RECT 63.920 152.225 64.330 152.555 ;
        RECT 61.450 151.795 62.300 151.965 ;
        RECT 62.860 151.575 63.180 152.035 ;
        RECT 63.380 151.785 63.630 152.215 ;
        RECT 63.920 151.575 64.330 152.015 ;
        RECT 64.500 151.955 64.670 152.685 ;
        RECT 64.840 152.135 65.190 152.505 ;
        RECT 65.370 152.195 65.590 153.065 ;
        RECT 65.760 152.495 66.170 153.115 ;
        RECT 66.340 152.315 66.510 153.285 ;
        RECT 65.815 152.125 66.510 152.315 ;
        RECT 64.500 151.755 65.515 151.955 ;
        RECT 65.815 151.795 65.985 152.125 ;
        RECT 66.155 151.575 66.485 151.955 ;
        RECT 66.700 151.835 66.925 153.955 ;
        RECT 67.095 153.625 67.425 154.125 ;
        RECT 67.595 153.455 67.765 153.955 ;
        RECT 67.100 153.285 67.765 153.455 ;
        RECT 67.100 152.295 67.330 153.285 ;
        RECT 67.500 152.465 67.850 153.115 ;
        RECT 68.485 153.035 71.075 154.125 ;
        RECT 71.335 153.195 71.505 153.955 ;
        RECT 71.720 153.365 72.050 154.125 ;
        RECT 68.485 152.515 69.695 153.035 ;
        RECT 71.335 153.025 72.050 153.195 ;
        RECT 72.220 153.050 72.475 153.955 ;
        RECT 69.865 152.345 71.075 152.865 ;
        RECT 71.245 152.475 71.600 152.845 ;
        RECT 71.880 152.815 72.050 153.025 ;
        RECT 71.880 152.485 72.135 152.815 ;
        RECT 67.100 152.125 67.765 152.295 ;
        RECT 67.095 151.575 67.425 151.955 ;
        RECT 67.595 151.835 67.765 152.125 ;
        RECT 68.485 151.575 71.075 152.345 ;
        RECT 71.880 152.295 72.050 152.485 ;
        RECT 72.305 152.320 72.475 153.050 ;
        RECT 72.650 152.975 72.910 154.125 ;
        RECT 73.095 153.065 73.425 154.125 ;
        RECT 73.605 152.815 73.775 153.785 ;
        RECT 73.945 153.535 74.275 153.935 ;
        RECT 74.445 153.765 74.775 154.125 ;
        RECT 74.975 153.535 75.675 153.955 ;
        RECT 73.945 153.305 75.675 153.535 ;
        RECT 73.945 153.085 74.275 153.305 ;
        RECT 74.470 152.815 74.795 153.105 ;
        RECT 73.085 152.485 73.395 152.815 ;
        RECT 73.605 152.485 73.980 152.815 ;
        RECT 74.300 152.485 74.795 152.815 ;
        RECT 74.970 152.565 75.300 153.105 ;
        RECT 71.335 152.125 72.050 152.295 ;
        RECT 71.335 151.745 71.505 152.125 ;
        RECT 71.720 151.575 72.050 151.955 ;
        RECT 72.220 151.745 72.475 152.320 ;
        RECT 72.650 151.575 72.910 152.415 ;
        RECT 75.470 152.335 75.675 153.305 ;
        RECT 75.845 152.960 76.135 154.125 ;
        RECT 77.225 153.035 80.735 154.125 ;
        RECT 80.910 153.690 86.255 154.125 ;
        RECT 77.225 152.515 78.915 153.035 ;
        RECT 79.085 152.345 80.735 152.865 ;
        RECT 82.500 152.440 82.850 153.690 ;
        RECT 86.800 153.145 87.055 153.815 ;
        RECT 87.235 153.325 87.520 154.125 ;
        RECT 87.700 153.405 88.030 153.915 ;
        RECT 73.095 152.105 74.455 152.315 ;
        RECT 73.095 151.745 73.425 152.105 ;
        RECT 73.595 151.575 73.925 151.935 ;
        RECT 74.125 151.745 74.455 152.105 ;
        RECT 74.965 151.745 75.675 152.335 ;
        RECT 75.845 151.575 76.135 152.300 ;
        RECT 77.225 151.575 80.735 152.345 ;
        RECT 84.330 152.120 84.670 152.950 ;
        RECT 86.800 152.285 86.980 153.145 ;
        RECT 87.700 152.815 87.950 153.405 ;
        RECT 88.300 153.255 88.470 153.865 ;
        RECT 88.640 153.435 88.970 154.125 ;
        RECT 89.200 153.575 89.440 153.865 ;
        RECT 89.640 153.745 90.060 154.125 ;
        RECT 90.240 153.655 90.870 153.905 ;
        RECT 91.340 153.745 91.670 154.125 ;
        RECT 90.240 153.575 90.410 153.655 ;
        RECT 91.840 153.575 92.010 153.865 ;
        RECT 92.190 153.745 92.570 154.125 ;
        RECT 92.810 153.740 93.640 153.910 ;
        RECT 89.200 153.405 90.410 153.575 ;
        RECT 87.150 152.485 87.950 152.815 ;
        RECT 80.910 151.575 86.255 152.120 ;
        RECT 86.800 152.085 87.055 152.285 ;
        RECT 86.715 151.915 87.055 152.085 ;
        RECT 86.800 151.755 87.055 151.915 ;
        RECT 87.235 151.575 87.520 152.035 ;
        RECT 87.700 151.835 87.950 152.485 ;
        RECT 88.150 153.235 88.470 153.255 ;
        RECT 88.150 153.065 90.070 153.235 ;
        RECT 88.150 152.170 88.340 153.065 ;
        RECT 90.240 152.895 90.410 153.405 ;
        RECT 90.580 153.145 91.100 153.455 ;
        RECT 88.510 152.725 90.410 152.895 ;
        RECT 88.510 152.665 88.840 152.725 ;
        RECT 88.990 152.495 89.320 152.555 ;
        RECT 88.660 152.225 89.320 152.495 ;
        RECT 88.150 151.840 88.470 152.170 ;
        RECT 88.650 151.575 89.310 152.055 ;
        RECT 89.510 151.965 89.680 152.725 ;
        RECT 90.580 152.555 90.760 152.965 ;
        RECT 89.850 152.385 90.180 152.505 ;
        RECT 90.930 152.385 91.100 153.145 ;
        RECT 89.850 152.215 91.100 152.385 ;
        RECT 91.270 153.325 92.640 153.575 ;
        RECT 91.270 152.555 91.460 153.325 ;
        RECT 92.390 153.065 92.640 153.325 ;
        RECT 91.630 152.895 91.880 153.055 ;
        RECT 92.810 152.895 92.980 153.740 ;
        RECT 93.875 153.455 94.045 153.955 ;
        RECT 94.215 153.625 94.545 154.125 ;
        RECT 93.150 153.065 93.650 153.445 ;
        RECT 93.875 153.285 94.570 153.455 ;
        RECT 91.630 152.725 92.980 152.895 ;
        RECT 92.560 152.685 92.980 152.725 ;
        RECT 91.270 152.215 91.690 152.555 ;
        RECT 91.980 152.225 92.390 152.555 ;
        RECT 89.510 151.795 90.360 151.965 ;
        RECT 90.920 151.575 91.240 152.035 ;
        RECT 91.440 151.785 91.690 152.215 ;
        RECT 91.980 151.575 92.390 152.015 ;
        RECT 92.560 151.955 92.730 152.685 ;
        RECT 92.900 152.135 93.250 152.505 ;
        RECT 93.430 152.195 93.650 153.065 ;
        RECT 93.820 152.495 94.230 153.115 ;
        RECT 94.400 152.315 94.570 153.285 ;
        RECT 93.875 152.125 94.570 152.315 ;
        RECT 92.560 151.755 93.575 151.955 ;
        RECT 93.875 151.795 94.045 152.125 ;
        RECT 94.215 151.575 94.545 151.955 ;
        RECT 94.760 151.835 94.985 153.955 ;
        RECT 95.155 153.625 95.485 154.125 ;
        RECT 95.655 153.455 95.825 153.955 ;
        RECT 96.090 153.690 101.435 154.125 ;
        RECT 95.160 153.285 95.825 153.455 ;
        RECT 95.160 152.295 95.390 153.285 ;
        RECT 95.560 152.465 95.910 153.115 ;
        RECT 97.680 152.440 98.030 153.690 ;
        RECT 101.605 152.960 101.895 154.125 ;
        RECT 102.525 152.985 102.795 153.955 ;
        RECT 103.005 153.325 103.285 154.125 ;
        RECT 103.455 153.615 105.110 153.905 ;
        RECT 103.520 153.275 105.110 153.445 ;
        RECT 103.520 153.155 103.690 153.275 ;
        RECT 102.965 152.985 103.690 153.155 ;
        RECT 95.160 152.125 95.825 152.295 ;
        RECT 95.155 151.575 95.485 151.955 ;
        RECT 95.655 151.835 95.825 152.125 ;
        RECT 99.510 152.120 99.850 152.950 ;
        RECT 96.090 151.575 101.435 152.120 ;
        RECT 101.605 151.575 101.895 152.300 ;
        RECT 102.525 152.250 102.695 152.985 ;
        RECT 102.965 152.815 103.135 152.985 ;
        RECT 103.880 152.935 104.595 153.105 ;
        RECT 104.790 152.985 105.110 153.275 ;
        RECT 105.285 152.985 105.625 153.955 ;
        RECT 105.795 152.985 105.965 154.125 ;
        RECT 106.235 153.325 106.485 154.125 ;
        RECT 107.130 153.155 107.460 153.955 ;
        RECT 107.760 153.325 108.090 154.125 ;
        RECT 108.260 153.155 108.590 153.955 ;
        RECT 106.155 152.985 108.590 153.155 ;
        RECT 108.965 152.985 109.305 153.955 ;
        RECT 109.475 152.985 109.645 154.125 ;
        RECT 109.915 153.325 110.165 154.125 ;
        RECT 110.810 153.155 111.140 153.955 ;
        RECT 111.440 153.325 111.770 154.125 ;
        RECT 111.940 153.155 112.270 153.955 ;
        RECT 113.110 153.690 118.455 154.125 ;
        RECT 109.835 152.985 112.270 153.155 ;
        RECT 102.865 152.485 103.135 152.815 ;
        RECT 103.305 152.485 103.710 152.815 ;
        RECT 103.880 152.485 104.590 152.935 ;
        RECT 102.965 152.315 103.135 152.485 ;
        RECT 102.525 151.905 102.795 152.250 ;
        RECT 102.965 152.145 104.575 152.315 ;
        RECT 104.760 152.245 105.110 152.815 ;
        RECT 105.285 152.375 105.460 152.985 ;
        RECT 106.155 152.735 106.325 152.985 ;
        RECT 105.630 152.565 106.325 152.735 ;
        RECT 106.500 152.565 106.920 152.765 ;
        RECT 107.090 152.565 107.420 152.765 ;
        RECT 107.590 152.565 107.920 152.765 ;
        RECT 102.985 151.575 103.365 151.975 ;
        RECT 103.535 151.795 103.705 152.145 ;
        RECT 103.875 151.575 104.205 151.975 ;
        RECT 104.405 151.795 104.575 152.145 ;
        RECT 104.775 151.575 105.105 152.075 ;
        RECT 105.285 151.745 105.625 152.375 ;
        RECT 105.795 151.575 106.045 152.375 ;
        RECT 106.235 152.225 107.460 152.395 ;
        RECT 106.235 151.745 106.565 152.225 ;
        RECT 106.735 151.575 106.960 152.035 ;
        RECT 107.130 151.745 107.460 152.225 ;
        RECT 108.090 152.355 108.260 152.985 ;
        RECT 108.445 152.565 108.795 152.815 ;
        RECT 108.965 152.425 109.140 152.985 ;
        RECT 109.835 152.735 110.005 152.985 ;
        RECT 109.310 152.565 110.005 152.735 ;
        RECT 110.180 152.565 110.600 152.765 ;
        RECT 110.770 152.565 111.100 152.765 ;
        RECT 111.270 152.565 111.600 152.765 ;
        RECT 108.965 152.375 109.195 152.425 ;
        RECT 108.090 151.745 108.590 152.355 ;
        RECT 108.965 151.745 109.305 152.375 ;
        RECT 109.475 151.575 109.725 152.375 ;
        RECT 109.915 152.225 111.140 152.395 ;
        RECT 109.915 151.745 110.245 152.225 ;
        RECT 110.415 151.575 110.640 152.035 ;
        RECT 110.810 151.745 111.140 152.225 ;
        RECT 111.770 152.355 111.940 152.985 ;
        RECT 112.125 152.565 112.475 152.815 ;
        RECT 114.700 152.440 115.050 153.690 ;
        RECT 118.685 152.985 118.895 154.125 ;
        RECT 119.065 152.975 119.395 153.955 ;
        RECT 119.565 152.985 119.795 154.125 ;
        RECT 120.555 153.195 120.725 153.955 ;
        RECT 120.905 153.365 121.235 154.125 ;
        RECT 120.555 153.025 121.220 153.195 ;
        RECT 121.405 153.050 121.675 153.955 ;
        RECT 111.770 151.745 112.270 152.355 ;
        RECT 116.530 152.120 116.870 152.950 ;
        RECT 113.110 151.575 118.455 152.120 ;
        RECT 118.685 151.575 118.895 152.395 ;
        RECT 119.065 152.375 119.315 152.975 ;
        RECT 121.050 152.880 121.220 153.025 ;
        RECT 119.485 152.565 119.815 152.815 ;
        RECT 120.485 152.475 120.815 152.845 ;
        RECT 121.050 152.550 121.335 152.880 ;
        RECT 119.065 151.745 119.395 152.375 ;
        RECT 119.565 151.575 119.795 152.395 ;
        RECT 121.050 152.295 121.220 152.550 ;
        RECT 120.555 152.125 121.220 152.295 ;
        RECT 121.505 152.250 121.675 153.050 ;
        RECT 122.765 153.035 126.275 154.125 ;
        RECT 126.445 153.035 127.655 154.125 ;
        RECT 122.765 152.515 124.455 153.035 ;
        RECT 124.625 152.345 126.275 152.865 ;
        RECT 126.445 152.495 126.965 153.035 ;
        RECT 120.555 151.745 120.725 152.125 ;
        RECT 120.905 151.575 121.235 151.955 ;
        RECT 121.415 151.745 121.675 152.250 ;
        RECT 122.765 151.575 126.275 152.345 ;
        RECT 127.135 152.325 127.655 152.865 ;
        RECT 126.445 151.575 127.655 152.325 ;
        RECT 14.580 151.405 127.740 151.575 ;
        RECT 14.665 150.655 15.875 151.405 ;
        RECT 16.880 150.695 17.135 151.225 ;
        RECT 17.315 150.945 17.600 151.405 ;
        RECT 14.665 150.115 15.185 150.655 ;
        RECT 15.355 149.945 15.875 150.485 ;
        RECT 16.880 150.045 17.060 150.695 ;
        RECT 17.780 150.495 18.030 151.145 ;
        RECT 17.230 150.165 18.030 150.495 ;
        RECT 14.665 148.855 15.875 149.945 ;
        RECT 16.795 149.875 17.060 150.045 ;
        RECT 16.880 149.835 17.060 149.875 ;
        RECT 16.880 149.165 17.135 149.835 ;
        RECT 17.315 148.855 17.600 149.655 ;
        RECT 17.780 149.575 18.030 150.165 ;
        RECT 18.230 150.810 18.550 151.140 ;
        RECT 18.730 150.925 19.390 151.405 ;
        RECT 19.590 151.015 20.440 151.185 ;
        RECT 18.230 149.915 18.420 150.810 ;
        RECT 18.740 150.485 19.400 150.755 ;
        RECT 19.070 150.425 19.400 150.485 ;
        RECT 18.590 150.255 18.920 150.315 ;
        RECT 19.590 150.255 19.760 151.015 ;
        RECT 21.000 150.945 21.320 151.405 ;
        RECT 21.520 150.765 21.770 151.195 ;
        RECT 22.060 150.965 22.470 151.405 ;
        RECT 22.640 151.025 23.655 151.225 ;
        RECT 19.930 150.595 21.180 150.765 ;
        RECT 19.930 150.475 20.260 150.595 ;
        RECT 18.590 150.085 20.490 150.255 ;
        RECT 18.230 149.745 20.150 149.915 ;
        RECT 18.230 149.725 18.550 149.745 ;
        RECT 17.780 149.065 18.110 149.575 ;
        RECT 18.380 149.115 18.550 149.725 ;
        RECT 20.320 149.575 20.490 150.085 ;
        RECT 20.660 150.015 20.840 150.425 ;
        RECT 21.010 149.835 21.180 150.595 ;
        RECT 18.720 148.855 19.050 149.545 ;
        RECT 19.280 149.405 20.490 149.575 ;
        RECT 20.660 149.525 21.180 149.835 ;
        RECT 21.350 150.425 21.770 150.765 ;
        RECT 22.060 150.425 22.470 150.755 ;
        RECT 21.350 149.655 21.540 150.425 ;
        RECT 22.640 150.295 22.810 151.025 ;
        RECT 23.955 150.855 24.125 151.185 ;
        RECT 24.295 151.025 24.625 151.405 ;
        RECT 22.980 150.475 23.330 150.845 ;
        RECT 22.640 150.255 23.060 150.295 ;
        RECT 21.710 150.085 23.060 150.255 ;
        RECT 21.710 149.925 21.960 150.085 ;
        RECT 22.470 149.655 22.720 149.915 ;
        RECT 21.350 149.405 22.720 149.655 ;
        RECT 19.280 149.115 19.520 149.405 ;
        RECT 20.320 149.325 20.490 149.405 ;
        RECT 19.720 148.855 20.140 149.235 ;
        RECT 20.320 149.075 20.950 149.325 ;
        RECT 21.420 148.855 21.750 149.235 ;
        RECT 21.920 149.115 22.090 149.405 ;
        RECT 22.890 149.240 23.060 150.085 ;
        RECT 23.510 149.915 23.730 150.785 ;
        RECT 23.955 150.665 24.650 150.855 ;
        RECT 23.230 149.535 23.730 149.915 ;
        RECT 23.900 149.865 24.310 150.485 ;
        RECT 24.480 149.695 24.650 150.665 ;
        RECT 23.955 149.525 24.650 149.695 ;
        RECT 22.270 148.855 22.650 149.235 ;
        RECT 22.890 149.070 23.720 149.240 ;
        RECT 23.955 149.025 24.125 149.525 ;
        RECT 24.295 148.855 24.625 149.355 ;
        RECT 24.840 149.025 25.065 151.145 ;
        RECT 25.235 151.025 25.565 151.405 ;
        RECT 25.735 150.855 25.905 151.145 ;
        RECT 25.240 150.685 25.905 150.855 ;
        RECT 25.240 149.695 25.470 150.685 ;
        RECT 26.165 150.655 27.375 151.405 ;
        RECT 27.550 150.860 32.895 151.405 ;
        RECT 25.640 149.865 25.990 150.515 ;
        RECT 26.165 149.945 26.685 150.485 ;
        RECT 26.855 150.115 27.375 150.655 ;
        RECT 25.240 149.525 25.905 149.695 ;
        RECT 25.235 148.855 25.565 149.355 ;
        RECT 25.735 149.025 25.905 149.525 ;
        RECT 26.165 148.855 27.375 149.945 ;
        RECT 29.140 149.290 29.490 150.540 ;
        RECT 30.970 150.030 31.310 150.860 ;
        RECT 33.105 150.585 33.335 151.405 ;
        RECT 33.505 150.605 33.835 151.235 ;
        RECT 33.085 150.165 33.415 150.415 ;
        RECT 33.585 150.005 33.835 150.605 ;
        RECT 34.005 150.585 34.215 151.405 ;
        RECT 34.445 150.655 35.655 151.405 ;
        RECT 35.915 150.855 36.085 151.235 ;
        RECT 36.265 151.025 36.595 151.405 ;
        RECT 35.915 150.685 36.580 150.855 ;
        RECT 36.775 150.730 37.035 151.235 ;
        RECT 27.550 148.855 32.895 149.290 ;
        RECT 33.105 148.855 33.335 149.995 ;
        RECT 33.505 149.025 33.835 150.005 ;
        RECT 34.005 148.855 34.215 149.995 ;
        RECT 34.445 149.945 34.965 150.485 ;
        RECT 35.135 150.115 35.655 150.655 ;
        RECT 35.845 150.135 36.175 150.505 ;
        RECT 36.410 150.430 36.580 150.685 ;
        RECT 36.410 150.100 36.695 150.430 ;
        RECT 36.410 149.955 36.580 150.100 ;
        RECT 34.445 148.855 35.655 149.945 ;
        RECT 35.915 149.785 36.580 149.955 ;
        RECT 36.865 149.930 37.035 150.730 ;
        RECT 37.205 150.680 37.495 151.405 ;
        RECT 37.665 150.635 41.175 151.405 ;
        RECT 35.915 149.025 36.085 149.785 ;
        RECT 36.265 148.855 36.595 149.615 ;
        RECT 36.765 149.025 37.035 149.930 ;
        RECT 37.205 148.855 37.495 150.020 ;
        RECT 37.665 149.945 39.355 150.465 ;
        RECT 39.525 150.115 41.175 150.635 ;
        RECT 41.345 150.605 41.685 151.235 ;
        RECT 41.855 150.605 42.105 151.405 ;
        RECT 42.295 150.755 42.625 151.235 ;
        RECT 42.795 150.945 43.020 151.405 ;
        RECT 43.190 150.755 43.520 151.235 ;
        RECT 41.345 149.995 41.520 150.605 ;
        RECT 42.295 150.585 43.520 150.755 ;
        RECT 44.150 150.625 44.650 151.235 ;
        RECT 45.025 150.635 48.535 151.405 ;
        RECT 48.715 150.905 49.045 151.405 ;
        RECT 49.245 150.835 49.415 151.185 ;
        RECT 49.615 151.005 49.945 151.405 ;
        RECT 50.115 150.835 50.285 151.185 ;
        RECT 50.455 151.005 50.835 151.405 ;
        RECT 41.690 150.245 42.385 150.415 ;
        RECT 42.215 149.995 42.385 150.245 ;
        RECT 42.560 150.215 42.980 150.415 ;
        RECT 43.150 150.215 43.480 150.415 ;
        RECT 43.650 150.215 43.980 150.415 ;
        RECT 44.150 149.995 44.320 150.625 ;
        RECT 44.505 150.165 44.855 150.415 ;
        RECT 37.665 148.855 41.175 149.945 ;
        RECT 41.345 149.025 41.685 149.995 ;
        RECT 41.855 148.855 42.025 149.995 ;
        RECT 42.215 149.825 44.650 149.995 ;
        RECT 42.295 148.855 42.545 149.655 ;
        RECT 43.190 149.025 43.520 149.825 ;
        RECT 43.820 148.855 44.150 149.655 ;
        RECT 44.320 149.025 44.650 149.825 ;
        RECT 45.025 149.945 46.715 150.465 ;
        RECT 46.885 150.115 48.535 150.635 ;
        RECT 48.710 150.165 49.060 150.735 ;
        RECT 49.245 150.665 50.855 150.835 ;
        RECT 51.025 150.730 51.295 151.075 ;
        RECT 50.685 150.495 50.855 150.665 ;
        RECT 45.025 148.855 48.535 149.945 ;
        RECT 48.710 149.705 49.030 149.995 ;
        RECT 49.230 149.875 49.940 150.495 ;
        RECT 50.110 150.165 50.515 150.495 ;
        RECT 50.685 150.165 50.955 150.495 ;
        RECT 50.685 149.995 50.855 150.165 ;
        RECT 51.125 149.995 51.295 150.730 ;
        RECT 50.130 149.825 50.855 149.995 ;
        RECT 50.130 149.705 50.300 149.825 ;
        RECT 48.710 149.535 50.300 149.705 ;
        RECT 48.710 149.075 50.365 149.365 ;
        RECT 50.535 148.855 50.815 149.655 ;
        RECT 51.025 149.025 51.295 149.995 ;
        RECT 51.465 150.605 51.805 151.235 ;
        RECT 51.975 150.605 52.225 151.405 ;
        RECT 52.415 150.755 52.745 151.235 ;
        RECT 52.915 150.945 53.140 151.405 ;
        RECT 53.310 150.755 53.640 151.235 ;
        RECT 51.465 149.995 51.640 150.605 ;
        RECT 52.415 150.585 53.640 150.755 ;
        RECT 54.270 150.625 54.770 151.235 ;
        RECT 55.145 150.635 56.815 151.405 ;
        RECT 51.810 150.245 52.505 150.415 ;
        RECT 52.335 149.995 52.505 150.245 ;
        RECT 52.680 150.215 53.100 150.415 ;
        RECT 53.270 150.215 53.600 150.415 ;
        RECT 53.770 150.215 54.100 150.415 ;
        RECT 54.270 149.995 54.440 150.625 ;
        RECT 54.625 150.165 54.975 150.415 ;
        RECT 51.465 149.025 51.805 149.995 ;
        RECT 51.975 148.855 52.145 149.995 ;
        RECT 52.335 149.825 54.770 149.995 ;
        RECT 52.415 148.855 52.665 149.655 ;
        RECT 53.310 149.025 53.640 149.825 ;
        RECT 53.940 148.855 54.270 149.655 ;
        RECT 54.440 149.025 54.770 149.825 ;
        RECT 55.145 149.945 55.895 150.465 ;
        RECT 56.065 150.115 56.815 150.635 ;
        RECT 57.260 150.595 57.505 151.200 ;
        RECT 57.725 150.870 58.235 151.405 ;
        RECT 56.985 150.425 58.215 150.595 ;
        RECT 55.145 148.855 56.815 149.945 ;
        RECT 56.985 149.615 57.325 150.425 ;
        RECT 57.495 149.860 58.245 150.050 ;
        RECT 56.985 149.205 57.500 149.615 ;
        RECT 57.735 148.855 57.905 149.615 ;
        RECT 58.075 149.195 58.245 149.860 ;
        RECT 58.415 149.875 58.605 151.235 ;
        RECT 58.775 150.385 59.050 151.235 ;
        RECT 59.240 150.870 59.770 151.235 ;
        RECT 60.195 151.005 60.525 151.405 ;
        RECT 59.595 150.835 59.770 150.870 ;
        RECT 58.775 150.215 59.055 150.385 ;
        RECT 58.775 150.075 59.050 150.215 ;
        RECT 59.255 149.875 59.425 150.675 ;
        RECT 58.415 149.705 59.425 149.875 ;
        RECT 59.595 150.665 60.525 150.835 ;
        RECT 60.695 150.665 60.950 151.235 ;
        RECT 59.595 149.535 59.765 150.665 ;
        RECT 60.355 150.495 60.525 150.665 ;
        RECT 58.640 149.365 59.765 149.535 ;
        RECT 59.935 150.165 60.130 150.495 ;
        RECT 60.355 150.165 60.610 150.495 ;
        RECT 59.935 149.195 60.105 150.165 ;
        RECT 60.780 149.995 60.950 150.665 ;
        RECT 58.075 149.025 60.105 149.195 ;
        RECT 60.275 148.855 60.445 149.995 ;
        RECT 60.615 149.025 60.950 149.995 ;
        RECT 61.585 150.730 61.845 151.235 ;
        RECT 62.025 151.025 62.355 151.405 ;
        RECT 62.535 150.855 62.705 151.235 ;
        RECT 61.585 149.930 61.755 150.730 ;
        RECT 62.040 150.685 62.705 150.855 ;
        RECT 62.040 150.430 62.210 150.685 ;
        RECT 62.965 150.680 63.255 151.405 ;
        RECT 63.975 150.855 64.145 151.235 ;
        RECT 64.325 151.025 64.655 151.405 ;
        RECT 63.975 150.685 64.640 150.855 ;
        RECT 64.835 150.730 65.095 151.235 ;
        RECT 61.925 150.100 62.210 150.430 ;
        RECT 62.445 150.135 62.775 150.505 ;
        RECT 63.905 150.135 64.235 150.505 ;
        RECT 64.470 150.430 64.640 150.685 ;
        RECT 62.040 149.955 62.210 150.100 ;
        RECT 64.470 150.100 64.755 150.430 ;
        RECT 61.585 149.025 61.855 149.930 ;
        RECT 62.040 149.785 62.705 149.955 ;
        RECT 62.025 148.855 62.355 149.615 ;
        RECT 62.535 149.025 62.705 149.785 ;
        RECT 62.965 148.855 63.255 150.020 ;
        RECT 64.470 149.955 64.640 150.100 ;
        RECT 63.975 149.785 64.640 149.955 ;
        RECT 64.925 149.930 65.095 150.730 ;
        RECT 65.725 150.635 67.395 151.405 ;
        RECT 67.655 150.855 67.825 151.235 ;
        RECT 68.040 151.025 68.370 151.405 ;
        RECT 67.655 150.685 68.370 150.855 ;
        RECT 63.975 149.025 64.145 149.785 ;
        RECT 64.325 148.855 64.655 149.615 ;
        RECT 64.825 149.025 65.095 149.930 ;
        RECT 65.725 149.945 66.475 150.465 ;
        RECT 66.645 150.115 67.395 150.635 ;
        RECT 67.565 150.135 67.920 150.505 ;
        RECT 68.200 150.495 68.370 150.685 ;
        RECT 68.540 150.660 68.795 151.235 ;
        RECT 68.200 150.165 68.455 150.495 ;
        RECT 68.200 149.955 68.370 150.165 ;
        RECT 65.725 148.855 67.395 149.945 ;
        RECT 67.655 149.785 68.370 149.955 ;
        RECT 68.625 149.930 68.795 150.660 ;
        RECT 68.970 150.565 69.230 151.405 ;
        RECT 69.410 150.565 69.670 151.405 ;
        RECT 69.845 150.660 70.100 151.235 ;
        RECT 70.270 151.025 70.600 151.405 ;
        RECT 70.815 150.855 70.985 151.235 ;
        RECT 71.305 150.925 71.585 151.405 ;
        RECT 70.270 150.685 70.985 150.855 ;
        RECT 71.755 150.755 72.015 151.145 ;
        RECT 72.190 150.925 72.445 151.405 ;
        RECT 72.615 150.755 72.910 151.145 ;
        RECT 73.090 150.925 73.365 151.405 ;
        RECT 73.535 150.905 73.835 151.235 ;
        RECT 67.655 149.025 67.825 149.785 ;
        RECT 68.040 148.855 68.370 149.615 ;
        RECT 68.540 149.025 68.795 149.930 ;
        RECT 68.970 148.855 69.230 150.005 ;
        RECT 69.410 148.855 69.670 150.005 ;
        RECT 69.845 149.930 70.015 150.660 ;
        RECT 70.270 150.495 70.440 150.685 ;
        RECT 71.260 150.585 72.910 150.755 ;
        RECT 70.185 150.165 70.440 150.495 ;
        RECT 70.270 149.955 70.440 150.165 ;
        RECT 70.720 150.135 71.075 150.505 ;
        RECT 71.260 150.075 71.665 150.585 ;
        RECT 71.835 150.245 72.975 150.415 ;
        RECT 69.845 149.025 70.100 149.930 ;
        RECT 70.270 149.785 70.985 149.955 ;
        RECT 71.260 149.905 72.015 150.075 ;
        RECT 70.270 148.855 70.600 149.615 ;
        RECT 70.815 149.025 70.985 149.785 ;
        RECT 71.300 148.855 71.585 149.725 ;
        RECT 71.755 149.655 72.015 149.905 ;
        RECT 72.805 149.995 72.975 150.245 ;
        RECT 73.145 150.165 73.495 150.735 ;
        RECT 73.665 149.995 73.835 150.905 ;
        RECT 72.805 149.825 73.835 149.995 ;
        RECT 71.755 149.485 72.875 149.655 ;
        RECT 71.755 149.025 72.015 149.485 ;
        RECT 72.190 148.855 72.445 149.315 ;
        RECT 72.615 149.025 72.875 149.485 ;
        RECT 73.045 148.855 73.355 149.655 ;
        RECT 73.525 149.025 73.835 149.825 ;
        RECT 74.925 150.905 75.225 151.235 ;
        RECT 75.395 150.925 75.670 151.405 ;
        RECT 74.925 149.995 75.095 150.905 ;
        RECT 75.850 150.755 76.145 151.145 ;
        RECT 76.315 150.925 76.570 151.405 ;
        RECT 76.745 150.755 77.005 151.145 ;
        RECT 77.175 150.925 77.455 151.405 ;
        RECT 75.265 150.165 75.615 150.735 ;
        RECT 75.850 150.585 77.500 150.755 ;
        RECT 75.785 150.245 76.925 150.415 ;
        RECT 75.785 149.995 75.955 150.245 ;
        RECT 77.095 150.075 77.500 150.585 ;
        RECT 74.925 149.825 75.955 149.995 ;
        RECT 76.745 149.905 77.500 150.075 ;
        RECT 77.685 150.730 77.955 151.075 ;
        RECT 78.145 151.005 78.525 151.405 ;
        RECT 78.695 150.835 78.865 151.185 ;
        RECT 79.035 151.005 79.365 151.405 ;
        RECT 79.565 150.835 79.735 151.185 ;
        RECT 79.935 150.905 80.265 151.405 ;
        RECT 77.685 149.995 77.855 150.730 ;
        RECT 78.125 150.665 79.735 150.835 ;
        RECT 78.125 150.495 78.295 150.665 ;
        RECT 78.025 150.165 78.295 150.495 ;
        RECT 78.465 150.165 78.870 150.495 ;
        RECT 78.125 149.995 78.295 150.165 ;
        RECT 79.040 150.045 79.750 150.495 ;
        RECT 79.920 150.165 80.270 150.735 ;
        RECT 80.905 150.635 84.415 151.405 ;
        RECT 74.925 149.025 75.235 149.825 ;
        RECT 76.745 149.655 77.005 149.905 ;
        RECT 75.405 148.855 75.715 149.655 ;
        RECT 75.885 149.485 77.005 149.655 ;
        RECT 75.885 149.025 76.145 149.485 ;
        RECT 76.315 148.855 76.570 149.315 ;
        RECT 76.745 149.025 77.005 149.485 ;
        RECT 77.175 148.855 77.460 149.725 ;
        RECT 77.685 149.025 77.955 149.995 ;
        RECT 78.125 149.825 78.850 149.995 ;
        RECT 79.040 149.875 79.755 150.045 ;
        RECT 78.680 149.705 78.850 149.825 ;
        RECT 79.950 149.705 80.270 149.995 ;
        RECT 78.165 148.855 78.445 149.655 ;
        RECT 78.680 149.535 80.270 149.705 ;
        RECT 80.905 149.945 82.595 150.465 ;
        RECT 82.765 150.115 84.415 150.635 ;
        RECT 84.860 150.595 85.105 151.200 ;
        RECT 85.325 150.870 85.835 151.405 ;
        RECT 84.585 150.425 85.815 150.595 ;
        RECT 78.615 149.075 80.270 149.365 ;
        RECT 80.905 148.855 84.415 149.945 ;
        RECT 84.585 149.615 84.925 150.425 ;
        RECT 85.095 149.860 85.845 150.050 ;
        RECT 84.585 149.205 85.100 149.615 ;
        RECT 85.335 148.855 85.505 149.615 ;
        RECT 85.675 149.195 85.845 149.860 ;
        RECT 86.015 149.875 86.205 151.235 ;
        RECT 86.375 150.385 86.650 151.235 ;
        RECT 86.840 150.870 87.370 151.235 ;
        RECT 87.795 151.005 88.125 151.405 ;
        RECT 87.195 150.835 87.370 150.870 ;
        RECT 86.375 150.215 86.655 150.385 ;
        RECT 86.375 150.075 86.650 150.215 ;
        RECT 86.855 149.875 87.025 150.675 ;
        RECT 86.015 149.705 87.025 149.875 ;
        RECT 87.195 150.665 88.125 150.835 ;
        RECT 88.295 150.665 88.550 151.235 ;
        RECT 88.725 150.680 89.015 151.405 ;
        RECT 87.195 149.535 87.365 150.665 ;
        RECT 87.955 150.495 88.125 150.665 ;
        RECT 86.240 149.365 87.365 149.535 ;
        RECT 87.535 150.165 87.730 150.495 ;
        RECT 87.955 150.165 88.210 150.495 ;
        RECT 87.535 149.195 87.705 150.165 ;
        RECT 88.380 149.995 88.550 150.665 ;
        RECT 89.705 150.585 89.915 151.405 ;
        RECT 90.085 150.605 90.415 151.235 ;
        RECT 85.675 149.025 87.705 149.195 ;
        RECT 87.875 148.855 88.045 149.995 ;
        RECT 88.215 149.025 88.550 149.995 ;
        RECT 88.725 148.855 89.015 150.020 ;
        RECT 90.085 150.005 90.335 150.605 ;
        RECT 90.585 150.585 90.815 151.405 ;
        RECT 92.035 150.855 92.205 151.235 ;
        RECT 92.385 151.025 92.715 151.405 ;
        RECT 92.035 150.685 92.700 150.855 ;
        RECT 92.895 150.730 93.155 151.235 ;
        RECT 90.505 150.165 90.835 150.415 ;
        RECT 91.965 150.135 92.295 150.505 ;
        RECT 92.530 150.430 92.700 150.685 ;
        RECT 92.530 150.100 92.815 150.430 ;
        RECT 89.705 148.855 89.915 149.995 ;
        RECT 90.085 149.025 90.415 150.005 ;
        RECT 90.585 148.855 90.815 149.995 ;
        RECT 92.530 149.955 92.700 150.100 ;
        RECT 92.035 149.785 92.700 149.955 ;
        RECT 92.985 149.930 93.155 150.730 ;
        RECT 93.385 150.585 93.595 151.405 ;
        RECT 93.765 150.605 94.095 151.235 ;
        RECT 93.765 150.005 94.015 150.605 ;
        RECT 94.265 150.585 94.495 151.405 ;
        RECT 94.705 150.635 96.375 151.405 ;
        RECT 94.185 150.165 94.515 150.415 ;
        RECT 92.035 149.025 92.205 149.785 ;
        RECT 92.385 148.855 92.715 149.615 ;
        RECT 92.885 149.025 93.155 149.930 ;
        RECT 93.385 148.855 93.595 149.995 ;
        RECT 93.765 149.025 94.095 150.005 ;
        RECT 94.265 148.855 94.495 149.995 ;
        RECT 94.705 149.945 95.455 150.465 ;
        RECT 95.625 150.115 96.375 150.635 ;
        RECT 96.550 150.695 96.805 151.225 ;
        RECT 96.975 150.945 97.280 151.405 ;
        RECT 97.525 151.025 98.595 151.195 ;
        RECT 96.550 150.045 96.760 150.695 ;
        RECT 97.525 150.670 97.845 151.025 ;
        RECT 97.520 150.495 97.845 150.670 ;
        RECT 96.930 150.195 97.845 150.495 ;
        RECT 98.015 150.455 98.255 150.855 ;
        RECT 98.425 150.795 98.595 151.025 ;
        RECT 98.765 150.965 98.955 151.405 ;
        RECT 99.125 150.955 100.075 151.235 ;
        RECT 100.295 151.045 100.645 151.215 ;
        RECT 98.425 150.625 98.955 150.795 ;
        RECT 96.930 150.165 97.670 150.195 ;
        RECT 94.705 148.855 96.375 149.945 ;
        RECT 96.550 149.165 96.805 150.045 ;
        RECT 96.975 148.855 97.280 149.995 ;
        RECT 97.500 149.575 97.670 150.165 ;
        RECT 98.015 150.085 98.555 150.455 ;
        RECT 98.735 150.345 98.955 150.625 ;
        RECT 99.125 150.175 99.295 150.955 ;
        RECT 98.890 150.005 99.295 150.175 ;
        RECT 99.465 150.165 99.815 150.785 ;
        RECT 98.890 149.915 99.060 150.005 ;
        RECT 99.985 149.995 100.195 150.785 ;
        RECT 97.840 149.745 99.060 149.915 ;
        RECT 99.520 149.835 100.195 149.995 ;
        RECT 97.500 149.405 98.300 149.575 ;
        RECT 97.620 148.855 97.950 149.235 ;
        RECT 98.130 149.115 98.300 149.405 ;
        RECT 98.890 149.365 99.060 149.745 ;
        RECT 99.230 149.825 100.195 149.835 ;
        RECT 100.385 150.655 100.645 151.045 ;
        RECT 100.855 150.945 101.185 151.405 ;
        RECT 102.060 151.015 102.915 151.185 ;
        RECT 103.120 151.015 103.615 151.185 ;
        RECT 103.785 151.045 104.115 151.405 ;
        RECT 100.385 149.965 100.555 150.655 ;
        RECT 100.725 150.305 100.895 150.485 ;
        RECT 101.065 150.475 101.855 150.725 ;
        RECT 102.060 150.305 102.230 151.015 ;
        RECT 102.400 150.505 102.755 150.725 ;
        RECT 100.725 150.135 102.415 150.305 ;
        RECT 99.230 149.535 99.690 149.825 ;
        RECT 100.385 149.795 101.885 149.965 ;
        RECT 100.385 149.655 100.555 149.795 ;
        RECT 99.995 149.485 100.555 149.655 ;
        RECT 98.470 148.855 98.720 149.315 ;
        RECT 98.890 149.025 99.760 149.365 ;
        RECT 99.995 149.025 100.165 149.485 ;
        RECT 101.000 149.455 102.075 149.625 ;
        RECT 100.335 148.855 100.705 149.315 ;
        RECT 101.000 149.115 101.170 149.455 ;
        RECT 101.340 148.855 101.670 149.285 ;
        RECT 101.905 149.115 102.075 149.455 ;
        RECT 102.245 149.355 102.415 150.135 ;
        RECT 102.585 149.915 102.755 150.505 ;
        RECT 102.925 150.105 103.275 150.725 ;
        RECT 102.585 149.525 103.050 149.915 ;
        RECT 103.445 149.655 103.615 151.015 ;
        RECT 103.785 149.825 104.245 150.875 ;
        RECT 103.220 149.485 103.615 149.655 ;
        RECT 103.220 149.355 103.390 149.485 ;
        RECT 102.245 149.025 102.925 149.355 ;
        RECT 103.140 149.025 103.390 149.355 ;
        RECT 103.560 148.855 103.810 149.315 ;
        RECT 103.980 149.040 104.305 149.825 ;
        RECT 104.475 149.025 104.645 151.145 ;
        RECT 104.815 151.025 105.145 151.405 ;
        RECT 105.315 150.855 105.570 151.145 ;
        RECT 104.820 150.685 105.570 150.855 ;
        RECT 104.820 149.695 105.050 150.685 ;
        RECT 105.745 150.655 106.955 151.405 ;
        RECT 105.220 149.865 105.570 150.515 ;
        RECT 105.745 149.945 106.265 150.485 ;
        RECT 106.435 150.115 106.955 150.655 ;
        RECT 107.125 150.605 107.465 151.235 ;
        RECT 107.635 150.605 107.885 151.405 ;
        RECT 108.075 150.755 108.405 151.235 ;
        RECT 108.575 150.945 108.800 151.405 ;
        RECT 108.970 150.755 109.300 151.235 ;
        RECT 107.125 149.995 107.300 150.605 ;
        RECT 108.075 150.585 109.300 150.755 ;
        RECT 109.930 150.625 110.430 151.235 ;
        RECT 110.920 150.775 111.205 151.235 ;
        RECT 111.375 150.945 111.645 151.405 ;
        RECT 107.470 150.245 108.165 150.415 ;
        RECT 107.995 149.995 108.165 150.245 ;
        RECT 108.340 150.215 108.760 150.415 ;
        RECT 108.930 150.215 109.260 150.415 ;
        RECT 109.430 150.215 109.760 150.415 ;
        RECT 109.930 149.995 110.100 150.625 ;
        RECT 110.920 150.605 111.875 150.775 ;
        RECT 110.285 150.165 110.635 150.415 ;
        RECT 104.820 149.525 105.570 149.695 ;
        RECT 104.815 148.855 105.145 149.355 ;
        RECT 105.315 149.025 105.570 149.525 ;
        RECT 105.745 148.855 106.955 149.945 ;
        RECT 107.125 149.025 107.465 149.995 ;
        RECT 107.635 148.855 107.805 149.995 ;
        RECT 107.995 149.825 110.430 149.995 ;
        RECT 110.805 149.875 111.495 150.435 ;
        RECT 108.075 148.855 108.325 149.655 ;
        RECT 108.970 149.025 109.300 149.825 ;
        RECT 109.600 148.855 109.930 149.655 ;
        RECT 110.100 149.025 110.430 149.825 ;
        RECT 111.665 149.705 111.875 150.605 ;
        RECT 110.920 149.485 111.875 149.705 ;
        RECT 112.045 150.435 112.445 151.235 ;
        RECT 112.635 150.775 112.915 151.235 ;
        RECT 113.435 150.945 113.760 151.405 ;
        RECT 112.635 150.605 113.760 150.775 ;
        RECT 113.930 150.665 114.315 151.235 ;
        RECT 114.485 150.680 114.775 151.405 ;
        RECT 115.870 150.695 116.125 151.225 ;
        RECT 116.295 150.945 116.600 151.405 ;
        RECT 116.845 151.025 117.915 151.195 ;
        RECT 113.310 150.495 113.760 150.605 ;
        RECT 112.045 149.875 113.140 150.435 ;
        RECT 113.310 150.165 113.865 150.495 ;
        RECT 110.920 149.025 111.205 149.485 ;
        RECT 111.375 148.855 111.645 149.315 ;
        RECT 112.045 149.025 112.445 149.875 ;
        RECT 113.310 149.705 113.760 150.165 ;
        RECT 114.035 149.995 114.315 150.665 ;
        RECT 115.870 150.045 116.080 150.695 ;
        RECT 116.845 150.670 117.165 151.025 ;
        RECT 116.840 150.495 117.165 150.670 ;
        RECT 116.250 150.195 117.165 150.495 ;
        RECT 117.335 150.455 117.575 150.855 ;
        RECT 117.745 150.795 117.915 151.025 ;
        RECT 118.085 150.965 118.275 151.405 ;
        RECT 118.445 150.955 119.395 151.235 ;
        RECT 119.615 151.045 119.965 151.215 ;
        RECT 117.745 150.625 118.275 150.795 ;
        RECT 116.250 150.165 116.990 150.195 ;
        RECT 112.635 149.485 113.760 149.705 ;
        RECT 112.635 149.025 112.915 149.485 ;
        RECT 113.435 148.855 113.760 149.315 ;
        RECT 113.930 149.025 114.315 149.995 ;
        RECT 114.485 148.855 114.775 150.020 ;
        RECT 115.870 149.165 116.125 150.045 ;
        RECT 116.295 148.855 116.600 149.995 ;
        RECT 116.820 149.575 116.990 150.165 ;
        RECT 117.335 150.085 117.875 150.455 ;
        RECT 118.055 150.345 118.275 150.625 ;
        RECT 118.445 150.175 118.615 150.955 ;
        RECT 118.210 150.005 118.615 150.175 ;
        RECT 118.785 150.165 119.135 150.785 ;
        RECT 118.210 149.915 118.380 150.005 ;
        RECT 119.305 149.995 119.515 150.785 ;
        RECT 117.160 149.745 118.380 149.915 ;
        RECT 118.840 149.835 119.515 149.995 ;
        RECT 116.820 149.405 117.620 149.575 ;
        RECT 116.940 148.855 117.270 149.235 ;
        RECT 117.450 149.115 117.620 149.405 ;
        RECT 118.210 149.365 118.380 149.745 ;
        RECT 118.550 149.825 119.515 149.835 ;
        RECT 119.705 150.655 119.965 151.045 ;
        RECT 120.175 150.945 120.505 151.405 ;
        RECT 121.380 151.015 122.235 151.185 ;
        RECT 122.440 151.015 122.935 151.185 ;
        RECT 123.105 151.045 123.435 151.405 ;
        RECT 119.705 149.965 119.875 150.655 ;
        RECT 120.045 150.305 120.215 150.485 ;
        RECT 120.385 150.475 121.175 150.725 ;
        RECT 121.380 150.305 121.550 151.015 ;
        RECT 121.720 150.505 122.075 150.725 ;
        RECT 120.045 150.135 121.735 150.305 ;
        RECT 118.550 149.535 119.010 149.825 ;
        RECT 119.705 149.795 121.205 149.965 ;
        RECT 119.705 149.655 119.875 149.795 ;
        RECT 119.315 149.485 119.875 149.655 ;
        RECT 117.790 148.855 118.040 149.315 ;
        RECT 118.210 149.025 119.080 149.365 ;
        RECT 119.315 149.025 119.485 149.485 ;
        RECT 120.320 149.455 121.395 149.625 ;
        RECT 119.655 148.855 120.025 149.315 ;
        RECT 120.320 149.115 120.490 149.455 ;
        RECT 120.660 148.855 120.990 149.285 ;
        RECT 121.225 149.115 121.395 149.455 ;
        RECT 121.565 149.355 121.735 150.135 ;
        RECT 121.905 149.915 122.075 150.505 ;
        RECT 122.245 150.105 122.595 150.725 ;
        RECT 121.905 149.525 122.370 149.915 ;
        RECT 122.765 149.655 122.935 151.015 ;
        RECT 123.105 149.825 123.565 150.875 ;
        RECT 122.540 149.485 122.935 149.655 ;
        RECT 122.540 149.355 122.710 149.485 ;
        RECT 121.565 149.025 122.245 149.355 ;
        RECT 122.460 149.025 122.710 149.355 ;
        RECT 122.880 148.855 123.130 149.315 ;
        RECT 123.300 149.040 123.625 149.825 ;
        RECT 123.795 149.025 123.965 151.145 ;
        RECT 124.135 151.025 124.465 151.405 ;
        RECT 124.635 150.855 124.890 151.145 ;
        RECT 124.140 150.685 124.890 150.855 ;
        RECT 124.140 149.695 124.370 150.685 ;
        RECT 125.065 150.655 126.275 151.405 ;
        RECT 126.445 150.655 127.655 151.405 ;
        RECT 124.540 149.865 124.890 150.515 ;
        RECT 125.065 149.945 125.585 150.485 ;
        RECT 125.755 150.115 126.275 150.655 ;
        RECT 126.445 149.945 126.965 150.485 ;
        RECT 127.135 150.115 127.655 150.655 ;
        RECT 124.140 149.525 124.890 149.695 ;
        RECT 124.135 148.855 124.465 149.355 ;
        RECT 124.635 149.025 124.890 149.525 ;
        RECT 125.065 148.855 126.275 149.945 ;
        RECT 126.445 148.855 127.655 149.945 ;
        RECT 14.580 148.685 127.740 148.855 ;
        RECT 14.665 147.595 15.875 148.685 ;
        RECT 14.665 146.885 15.185 147.425 ;
        RECT 15.355 147.055 15.875 147.595 ;
        RECT 16.505 147.595 20.015 148.685 ;
        RECT 20.185 147.925 20.700 148.335 ;
        RECT 20.935 147.925 21.105 148.685 ;
        RECT 21.275 148.345 23.305 148.515 ;
        RECT 16.505 147.075 18.195 147.595 ;
        RECT 18.365 146.905 20.015 147.425 ;
        RECT 20.185 147.115 20.525 147.925 ;
        RECT 21.275 147.680 21.445 148.345 ;
        RECT 21.840 148.005 22.965 148.175 ;
        RECT 20.695 147.490 21.445 147.680 ;
        RECT 21.615 147.665 22.625 147.835 ;
        RECT 20.185 146.945 21.415 147.115 ;
        RECT 14.665 146.135 15.875 146.885 ;
        RECT 16.505 146.135 20.015 146.905 ;
        RECT 20.460 146.340 20.705 146.945 ;
        RECT 20.925 146.135 21.435 146.670 ;
        RECT 21.615 146.305 21.805 147.665 ;
        RECT 21.975 146.985 22.250 147.465 ;
        RECT 21.975 146.815 22.255 146.985 ;
        RECT 22.455 146.865 22.625 147.665 ;
        RECT 22.795 146.875 22.965 148.005 ;
        RECT 23.135 147.375 23.305 148.345 ;
        RECT 23.475 147.545 23.645 148.685 ;
        RECT 23.815 147.545 24.150 148.515 ;
        RECT 23.135 147.045 23.330 147.375 ;
        RECT 23.555 147.045 23.810 147.375 ;
        RECT 23.555 146.875 23.725 147.045 ;
        RECT 23.980 146.875 24.150 147.545 ;
        RECT 24.325 147.520 24.615 148.685 ;
        RECT 24.785 147.610 25.055 148.515 ;
        RECT 25.225 147.925 25.555 148.685 ;
        RECT 25.735 147.755 25.905 148.515 ;
        RECT 21.975 146.305 22.250 146.815 ;
        RECT 22.795 146.705 23.725 146.875 ;
        RECT 22.795 146.670 22.970 146.705 ;
        RECT 22.440 146.305 22.970 146.670 ;
        RECT 23.395 146.135 23.725 146.535 ;
        RECT 23.895 146.305 24.150 146.875 ;
        RECT 24.325 146.135 24.615 146.860 ;
        RECT 24.785 146.810 24.955 147.610 ;
        RECT 25.240 147.585 25.905 147.755 ;
        RECT 26.165 147.595 27.835 148.685 ;
        RECT 28.095 147.755 28.265 148.515 ;
        RECT 28.445 147.925 28.775 148.685 ;
        RECT 25.240 147.440 25.410 147.585 ;
        RECT 25.125 147.110 25.410 147.440 ;
        RECT 25.240 146.855 25.410 147.110 ;
        RECT 25.645 147.035 25.975 147.405 ;
        RECT 26.165 147.075 26.915 147.595 ;
        RECT 28.095 147.585 28.760 147.755 ;
        RECT 28.945 147.610 29.215 148.515 ;
        RECT 28.590 147.440 28.760 147.585 ;
        RECT 27.085 146.905 27.835 147.425 ;
        RECT 28.025 147.035 28.355 147.405 ;
        RECT 28.590 147.110 28.875 147.440 ;
        RECT 24.785 146.305 25.045 146.810 ;
        RECT 25.240 146.685 25.905 146.855 ;
        RECT 25.225 146.135 25.555 146.515 ;
        RECT 25.735 146.305 25.905 146.685 ;
        RECT 26.165 146.135 27.835 146.905 ;
        RECT 28.590 146.855 28.760 147.110 ;
        RECT 28.095 146.685 28.760 146.855 ;
        RECT 29.045 146.810 29.215 147.610 ;
        RECT 28.095 146.305 28.265 146.685 ;
        RECT 28.445 146.135 28.775 146.515 ;
        RECT 28.955 146.305 29.215 146.810 ;
        RECT 29.390 147.545 29.725 148.515 ;
        RECT 29.895 147.545 30.065 148.685 ;
        RECT 30.235 148.345 32.265 148.515 ;
        RECT 29.390 146.875 29.560 147.545 ;
        RECT 30.235 147.375 30.405 148.345 ;
        RECT 29.730 147.045 29.985 147.375 ;
        RECT 30.210 147.045 30.405 147.375 ;
        RECT 30.575 148.005 31.700 148.175 ;
        RECT 29.815 146.875 29.985 147.045 ;
        RECT 30.575 146.875 30.745 148.005 ;
        RECT 29.390 146.305 29.645 146.875 ;
        RECT 29.815 146.705 30.745 146.875 ;
        RECT 30.915 147.665 31.925 147.835 ;
        RECT 30.915 146.865 31.085 147.665 ;
        RECT 31.290 147.325 31.565 147.465 ;
        RECT 31.285 147.155 31.565 147.325 ;
        RECT 30.570 146.670 30.745 146.705 ;
        RECT 29.815 146.135 30.145 146.535 ;
        RECT 30.570 146.305 31.100 146.670 ;
        RECT 31.290 146.305 31.565 147.155 ;
        RECT 31.735 146.305 31.925 147.665 ;
        RECT 32.095 147.680 32.265 148.345 ;
        RECT 32.435 147.925 32.605 148.685 ;
        RECT 32.840 147.925 33.355 148.335 ;
        RECT 32.095 147.490 32.845 147.680 ;
        RECT 33.015 147.115 33.355 147.925 ;
        RECT 32.125 146.945 33.355 147.115 ;
        RECT 33.985 147.595 35.655 148.685 ;
        RECT 36.030 147.715 36.360 148.515 ;
        RECT 36.530 147.885 36.860 148.685 ;
        RECT 37.160 147.715 37.490 148.515 ;
        RECT 38.135 147.885 38.385 148.685 ;
        RECT 33.985 147.075 34.735 147.595 ;
        RECT 36.030 147.545 38.465 147.715 ;
        RECT 38.655 147.545 38.825 148.685 ;
        RECT 38.995 147.545 39.335 148.515 ;
        RECT 32.105 146.135 32.615 146.670 ;
        RECT 32.835 146.340 33.080 146.945 ;
        RECT 34.905 146.905 35.655 147.425 ;
        RECT 35.825 147.125 36.175 147.375 ;
        RECT 36.360 146.915 36.530 147.545 ;
        RECT 36.700 147.125 37.030 147.325 ;
        RECT 37.200 147.125 37.530 147.325 ;
        RECT 37.700 147.125 38.120 147.325 ;
        RECT 38.295 147.295 38.465 147.545 ;
        RECT 38.295 147.125 38.990 147.295 ;
        RECT 33.985 146.135 35.655 146.905 ;
        RECT 36.030 146.305 36.530 146.915 ;
        RECT 37.160 146.785 38.385 146.955 ;
        RECT 39.160 146.935 39.335 147.545 ;
        RECT 37.160 146.305 37.490 146.785 ;
        RECT 37.660 146.135 37.885 146.595 ;
        RECT 38.055 146.305 38.385 146.785 ;
        RECT 38.575 146.135 38.825 146.935 ;
        RECT 38.995 146.305 39.335 146.935 ;
        RECT 39.505 147.545 39.845 148.515 ;
        RECT 40.015 147.545 40.185 148.685 ;
        RECT 40.455 147.885 40.705 148.685 ;
        RECT 41.350 147.715 41.680 148.515 ;
        RECT 41.980 147.885 42.310 148.685 ;
        RECT 42.480 147.715 42.810 148.515 ;
        RECT 40.375 147.545 42.810 147.715 ;
        RECT 43.645 147.595 47.155 148.685 ;
        RECT 47.330 148.175 48.985 148.465 ;
        RECT 47.330 147.835 48.920 148.005 ;
        RECT 49.155 147.885 49.435 148.685 ;
        RECT 39.505 146.985 39.680 147.545 ;
        RECT 40.375 147.295 40.545 147.545 ;
        RECT 39.850 147.125 40.545 147.295 ;
        RECT 40.720 147.125 41.140 147.325 ;
        RECT 41.310 147.125 41.640 147.325 ;
        RECT 41.810 147.125 42.140 147.325 ;
        RECT 39.505 146.935 39.735 146.985 ;
        RECT 39.505 146.305 39.845 146.935 ;
        RECT 40.015 146.135 40.265 146.935 ;
        RECT 40.455 146.785 41.680 146.955 ;
        RECT 40.455 146.305 40.785 146.785 ;
        RECT 40.955 146.135 41.180 146.595 ;
        RECT 41.350 146.305 41.680 146.785 ;
        RECT 42.310 146.915 42.480 147.545 ;
        RECT 42.665 147.125 43.015 147.375 ;
        RECT 43.645 147.075 45.335 147.595 ;
        RECT 47.330 147.545 47.650 147.835 ;
        RECT 48.750 147.715 48.920 147.835 ;
        RECT 42.310 146.305 42.810 146.915 ;
        RECT 45.505 146.905 47.155 147.425 ;
        RECT 43.645 146.135 47.155 146.905 ;
        RECT 47.330 146.805 47.680 147.375 ;
        RECT 47.850 147.045 48.560 147.665 ;
        RECT 48.750 147.545 49.475 147.715 ;
        RECT 49.645 147.545 49.915 148.515 ;
        RECT 49.305 147.375 49.475 147.545 ;
        RECT 48.730 147.045 49.135 147.375 ;
        RECT 49.305 147.045 49.575 147.375 ;
        RECT 49.305 146.875 49.475 147.045 ;
        RECT 47.865 146.705 49.475 146.875 ;
        RECT 49.745 146.810 49.915 147.545 ;
        RECT 50.085 147.520 50.375 148.685 ;
        RECT 51.005 147.610 51.275 148.515 ;
        RECT 51.445 147.925 51.775 148.685 ;
        RECT 51.955 147.755 52.125 148.515 ;
        RECT 47.335 146.135 47.665 146.635 ;
        RECT 47.865 146.355 48.035 146.705 ;
        RECT 48.235 146.135 48.565 146.535 ;
        RECT 48.735 146.355 48.905 146.705 ;
        RECT 49.075 146.135 49.455 146.535 ;
        RECT 49.645 146.465 49.915 146.810 ;
        RECT 50.085 146.135 50.375 146.860 ;
        RECT 51.005 146.810 51.175 147.610 ;
        RECT 51.460 147.585 52.125 147.755 ;
        RECT 51.460 147.440 51.630 147.585 ;
        RECT 51.345 147.110 51.630 147.440 ;
        RECT 53.305 147.545 53.645 148.515 ;
        RECT 53.815 147.545 53.985 148.685 ;
        RECT 54.255 147.885 54.505 148.685 ;
        RECT 55.150 147.715 55.480 148.515 ;
        RECT 55.780 147.885 56.110 148.685 ;
        RECT 56.280 147.715 56.610 148.515 ;
        RECT 54.175 147.545 56.610 147.715 ;
        RECT 56.985 147.595 59.575 148.685 ;
        RECT 59.745 147.925 60.260 148.335 ;
        RECT 60.495 147.925 60.665 148.685 ;
        RECT 60.835 148.345 62.865 148.515 ;
        RECT 51.460 146.855 51.630 147.110 ;
        RECT 51.865 147.035 52.195 147.405 ;
        RECT 53.305 146.935 53.480 147.545 ;
        RECT 54.175 147.295 54.345 147.545 ;
        RECT 53.650 147.125 54.345 147.295 ;
        RECT 54.520 147.125 54.940 147.325 ;
        RECT 55.110 147.125 55.440 147.325 ;
        RECT 55.610 147.125 55.940 147.325 ;
        RECT 51.005 146.305 51.265 146.810 ;
        RECT 51.460 146.685 52.125 146.855 ;
        RECT 51.445 146.135 51.775 146.515 ;
        RECT 51.955 146.305 52.125 146.685 ;
        RECT 53.305 146.305 53.645 146.935 ;
        RECT 53.815 146.135 54.065 146.935 ;
        RECT 54.255 146.785 55.480 146.955 ;
        RECT 54.255 146.305 54.585 146.785 ;
        RECT 54.755 146.135 54.980 146.595 ;
        RECT 55.150 146.305 55.480 146.785 ;
        RECT 56.110 146.915 56.280 147.545 ;
        RECT 56.465 147.125 56.815 147.375 ;
        RECT 56.985 147.075 58.195 147.595 ;
        RECT 56.110 146.305 56.610 146.915 ;
        RECT 58.365 146.905 59.575 147.425 ;
        RECT 59.745 147.115 60.085 147.925 ;
        RECT 60.835 147.680 61.005 148.345 ;
        RECT 61.400 148.005 62.525 148.175 ;
        RECT 60.255 147.490 61.005 147.680 ;
        RECT 61.175 147.665 62.185 147.835 ;
        RECT 59.745 146.945 60.975 147.115 ;
        RECT 56.985 146.135 59.575 146.905 ;
        RECT 60.020 146.340 60.265 146.945 ;
        RECT 60.485 146.135 60.995 146.670 ;
        RECT 61.175 146.305 61.365 147.665 ;
        RECT 61.535 146.645 61.810 147.465 ;
        RECT 62.015 146.865 62.185 147.665 ;
        RECT 62.355 146.875 62.525 148.005 ;
        RECT 62.695 147.375 62.865 148.345 ;
        RECT 63.035 147.545 63.205 148.685 ;
        RECT 63.375 147.545 63.710 148.515 ;
        RECT 62.695 147.045 62.890 147.375 ;
        RECT 63.115 147.045 63.370 147.375 ;
        RECT 63.115 146.875 63.285 147.045 ;
        RECT 63.540 146.875 63.710 147.545 ;
        RECT 63.885 147.595 65.095 148.685 ;
        RECT 65.270 148.250 70.615 148.685 ;
        RECT 63.885 147.055 64.405 147.595 ;
        RECT 64.575 146.885 65.095 147.425 ;
        RECT 66.860 147.000 67.210 148.250 ;
        RECT 70.790 147.535 71.050 148.685 ;
        RECT 71.225 147.610 71.480 148.515 ;
        RECT 71.650 147.925 71.980 148.685 ;
        RECT 72.195 147.755 72.365 148.515 ;
        RECT 62.355 146.705 63.285 146.875 ;
        RECT 62.355 146.670 62.530 146.705 ;
        RECT 61.535 146.475 61.815 146.645 ;
        RECT 61.535 146.305 61.810 146.475 ;
        RECT 62.000 146.305 62.530 146.670 ;
        RECT 62.955 146.135 63.285 146.535 ;
        RECT 63.455 146.305 63.710 146.875 ;
        RECT 63.885 146.135 65.095 146.885 ;
        RECT 68.690 146.680 69.030 147.510 ;
        RECT 65.270 146.135 70.615 146.680 ;
        RECT 70.790 146.135 71.050 146.975 ;
        RECT 71.225 146.880 71.395 147.610 ;
        RECT 71.650 147.585 72.365 147.755 ;
        RECT 72.715 147.755 72.885 148.515 ;
        RECT 73.100 147.925 73.430 148.685 ;
        RECT 72.715 147.585 73.430 147.755 ;
        RECT 73.600 147.610 73.855 148.515 ;
        RECT 71.650 147.375 71.820 147.585 ;
        RECT 71.565 147.045 71.820 147.375 ;
        RECT 71.225 146.305 71.480 146.880 ;
        RECT 71.650 146.855 71.820 147.045 ;
        RECT 72.100 147.035 72.455 147.405 ;
        RECT 72.625 147.035 72.980 147.405 ;
        RECT 73.260 147.375 73.430 147.585 ;
        RECT 73.260 147.045 73.515 147.375 ;
        RECT 73.260 146.855 73.430 147.045 ;
        RECT 73.685 146.880 73.855 147.610 ;
        RECT 74.030 147.535 74.290 148.685 ;
        RECT 74.465 147.595 75.675 148.685 ;
        RECT 74.465 147.055 74.985 147.595 ;
        RECT 75.845 147.520 76.135 148.685 ;
        RECT 76.510 147.715 76.840 148.515 ;
        RECT 77.010 147.885 77.340 148.685 ;
        RECT 77.640 147.715 77.970 148.515 ;
        RECT 78.615 147.885 78.865 148.685 ;
        RECT 76.510 147.545 78.945 147.715 ;
        RECT 79.135 147.545 79.305 148.685 ;
        RECT 79.475 147.545 79.815 148.515 ;
        RECT 71.650 146.685 72.365 146.855 ;
        RECT 71.650 146.135 71.980 146.515 ;
        RECT 72.195 146.305 72.365 146.685 ;
        RECT 72.715 146.685 73.430 146.855 ;
        RECT 72.715 146.305 72.885 146.685 ;
        RECT 73.100 146.135 73.430 146.515 ;
        RECT 73.600 146.305 73.855 146.880 ;
        RECT 74.030 146.135 74.290 146.975 ;
        RECT 75.155 146.885 75.675 147.425 ;
        RECT 76.305 147.125 76.655 147.375 ;
        RECT 76.840 146.915 77.010 147.545 ;
        RECT 77.180 147.125 77.510 147.325 ;
        RECT 77.680 147.125 78.010 147.325 ;
        RECT 78.180 147.125 78.600 147.325 ;
        RECT 78.775 147.295 78.945 147.545 ;
        RECT 78.775 147.125 79.470 147.295 ;
        RECT 74.465 146.135 75.675 146.885 ;
        RECT 75.845 146.135 76.135 146.860 ;
        RECT 76.510 146.305 77.010 146.915 ;
        RECT 77.640 146.785 78.865 146.955 ;
        RECT 79.640 146.935 79.815 147.545 ;
        RECT 77.640 146.305 77.970 146.785 ;
        RECT 78.140 146.135 78.365 146.595 ;
        RECT 78.535 146.305 78.865 146.785 ;
        RECT 79.055 146.135 79.305 146.935 ;
        RECT 79.475 146.305 79.815 146.935 ;
        RECT 79.985 147.545 80.325 148.515 ;
        RECT 80.495 147.545 80.665 148.685 ;
        RECT 80.935 147.885 81.185 148.685 ;
        RECT 81.830 147.715 82.160 148.515 ;
        RECT 82.460 147.885 82.790 148.685 ;
        RECT 82.960 147.715 83.290 148.515 ;
        RECT 80.855 147.545 83.290 147.715 ;
        RECT 83.665 147.595 84.875 148.685 ;
        RECT 85.420 147.705 85.675 148.375 ;
        RECT 85.855 147.885 86.140 148.685 ;
        RECT 86.320 147.965 86.650 148.475 ;
        RECT 79.985 146.935 80.160 147.545 ;
        RECT 80.855 147.295 81.025 147.545 ;
        RECT 80.330 147.125 81.025 147.295 ;
        RECT 81.200 147.125 81.620 147.325 ;
        RECT 81.790 147.125 82.120 147.325 ;
        RECT 82.290 147.125 82.620 147.325 ;
        RECT 79.985 146.305 80.325 146.935 ;
        RECT 80.495 146.135 80.745 146.935 ;
        RECT 80.935 146.785 82.160 146.955 ;
        RECT 80.935 146.305 81.265 146.785 ;
        RECT 81.435 146.135 81.660 146.595 ;
        RECT 81.830 146.305 82.160 146.785 ;
        RECT 82.790 146.915 82.960 147.545 ;
        RECT 83.145 147.125 83.495 147.375 ;
        RECT 83.665 147.055 84.185 147.595 ;
        RECT 82.790 146.305 83.290 146.915 ;
        RECT 84.355 146.885 84.875 147.425 ;
        RECT 83.665 146.135 84.875 146.885 ;
        RECT 85.420 146.845 85.600 147.705 ;
        RECT 86.320 147.375 86.570 147.965 ;
        RECT 86.920 147.815 87.090 148.425 ;
        RECT 87.260 147.995 87.590 148.685 ;
        RECT 87.820 148.135 88.060 148.425 ;
        RECT 88.260 148.305 88.680 148.685 ;
        RECT 88.860 148.215 89.490 148.465 ;
        RECT 89.960 148.305 90.290 148.685 ;
        RECT 88.860 148.135 89.030 148.215 ;
        RECT 90.460 148.135 90.630 148.425 ;
        RECT 90.810 148.305 91.190 148.685 ;
        RECT 91.430 148.300 92.260 148.470 ;
        RECT 87.820 147.965 89.030 148.135 ;
        RECT 85.770 147.045 86.570 147.375 ;
        RECT 85.420 146.645 85.675 146.845 ;
        RECT 85.335 146.475 85.675 146.645 ;
        RECT 85.420 146.315 85.675 146.475 ;
        RECT 85.855 146.135 86.140 146.595 ;
        RECT 86.320 146.395 86.570 147.045 ;
        RECT 86.770 147.795 87.090 147.815 ;
        RECT 86.770 147.625 88.690 147.795 ;
        RECT 86.770 146.730 86.960 147.625 ;
        RECT 88.860 147.455 89.030 147.965 ;
        RECT 89.200 147.705 89.720 148.015 ;
        RECT 87.130 147.285 89.030 147.455 ;
        RECT 87.130 147.225 87.460 147.285 ;
        RECT 87.610 147.055 87.940 147.115 ;
        RECT 87.280 146.785 87.940 147.055 ;
        RECT 86.770 146.400 87.090 146.730 ;
        RECT 87.270 146.135 87.930 146.615 ;
        RECT 88.130 146.525 88.300 147.285 ;
        RECT 89.200 147.115 89.380 147.525 ;
        RECT 88.470 146.945 88.800 147.065 ;
        RECT 89.550 146.945 89.720 147.705 ;
        RECT 88.470 146.775 89.720 146.945 ;
        RECT 89.890 147.885 91.260 148.135 ;
        RECT 89.890 147.115 90.080 147.885 ;
        RECT 91.010 147.625 91.260 147.885 ;
        RECT 90.250 147.455 90.500 147.615 ;
        RECT 91.430 147.455 91.600 148.300 ;
        RECT 92.495 148.015 92.665 148.515 ;
        RECT 92.835 148.185 93.165 148.685 ;
        RECT 91.770 147.625 92.270 148.005 ;
        RECT 92.495 147.845 93.190 148.015 ;
        RECT 90.250 147.285 91.600 147.455 ;
        RECT 91.180 147.245 91.600 147.285 ;
        RECT 89.890 146.775 90.310 147.115 ;
        RECT 90.600 146.785 91.010 147.115 ;
        RECT 88.130 146.355 88.980 146.525 ;
        RECT 89.540 146.135 89.860 146.595 ;
        RECT 90.060 146.345 90.310 146.775 ;
        RECT 90.600 146.135 91.010 146.575 ;
        RECT 91.180 146.515 91.350 147.245 ;
        RECT 91.520 146.695 91.870 147.065 ;
        RECT 92.050 146.755 92.270 147.625 ;
        RECT 92.440 147.055 92.850 147.675 ;
        RECT 93.020 146.875 93.190 147.845 ;
        RECT 92.495 146.685 93.190 146.875 ;
        RECT 91.180 146.315 92.195 146.515 ;
        RECT 92.495 146.355 92.665 146.685 ;
        RECT 92.835 146.135 93.165 146.515 ;
        RECT 93.380 146.395 93.605 148.515 ;
        RECT 93.775 148.185 94.105 148.685 ;
        RECT 94.275 148.015 94.445 148.515 ;
        RECT 93.780 147.845 94.445 148.015 ;
        RECT 93.780 146.855 94.010 147.845 ;
        RECT 94.180 147.025 94.530 147.675 ;
        RECT 95.205 147.545 95.435 148.685 ;
        RECT 95.605 147.535 95.935 148.515 ;
        RECT 96.105 147.545 96.315 148.685 ;
        RECT 96.545 147.925 97.060 148.335 ;
        RECT 97.295 147.925 97.465 148.685 ;
        RECT 97.635 148.345 99.665 148.515 ;
        RECT 95.185 147.125 95.515 147.375 ;
        RECT 93.780 146.685 94.445 146.855 ;
        RECT 93.775 146.135 94.105 146.515 ;
        RECT 94.275 146.395 94.445 146.685 ;
        RECT 95.205 146.135 95.435 146.955 ;
        RECT 95.685 146.935 95.935 147.535 ;
        RECT 96.545 147.115 96.885 147.925 ;
        RECT 97.635 147.680 97.805 148.345 ;
        RECT 98.200 148.005 99.325 148.175 ;
        RECT 97.055 147.490 97.805 147.680 ;
        RECT 97.975 147.665 98.985 147.835 ;
        RECT 95.605 146.305 95.935 146.935 ;
        RECT 96.105 146.135 96.315 146.955 ;
        RECT 96.545 146.945 97.775 147.115 ;
        RECT 96.820 146.340 97.065 146.945 ;
        RECT 97.285 146.135 97.795 146.670 ;
        RECT 97.975 146.305 98.165 147.665 ;
        RECT 98.335 147.325 98.610 147.465 ;
        RECT 98.335 147.155 98.615 147.325 ;
        RECT 98.335 146.305 98.610 147.155 ;
        RECT 98.815 146.865 98.985 147.665 ;
        RECT 99.155 146.875 99.325 148.005 ;
        RECT 99.495 147.375 99.665 148.345 ;
        RECT 99.835 147.545 100.005 148.685 ;
        RECT 100.175 147.545 100.510 148.515 ;
        RECT 99.495 147.045 99.690 147.375 ;
        RECT 99.915 147.045 100.170 147.375 ;
        RECT 99.915 146.875 100.085 147.045 ;
        RECT 100.340 146.875 100.510 147.545 ;
        RECT 101.605 147.520 101.895 148.685 ;
        RECT 102.155 147.755 102.325 148.515 ;
        RECT 102.505 147.925 102.835 148.685 ;
        RECT 102.155 147.585 102.820 147.755 ;
        RECT 103.005 147.610 103.275 148.515 ;
        RECT 102.650 147.440 102.820 147.585 ;
        RECT 102.085 147.035 102.415 147.405 ;
        RECT 102.650 147.110 102.935 147.440 ;
        RECT 99.155 146.705 100.085 146.875 ;
        RECT 99.155 146.670 99.330 146.705 ;
        RECT 98.800 146.305 99.330 146.670 ;
        RECT 99.755 146.135 100.085 146.535 ;
        RECT 100.255 146.305 100.510 146.875 ;
        RECT 101.605 146.135 101.895 146.860 ;
        RECT 102.650 146.855 102.820 147.110 ;
        RECT 102.155 146.685 102.820 146.855 ;
        RECT 103.105 146.810 103.275 147.610 ;
        RECT 102.155 146.305 102.325 146.685 ;
        RECT 102.505 146.135 102.835 146.515 ;
        RECT 103.015 146.305 103.275 146.810 ;
        RECT 103.905 147.545 104.175 148.515 ;
        RECT 104.385 147.885 104.665 148.685 ;
        RECT 104.835 148.175 106.490 148.465 ;
        RECT 104.900 147.835 106.490 148.005 ;
        RECT 104.900 147.715 105.070 147.835 ;
        RECT 104.345 147.545 105.070 147.715 ;
        RECT 103.905 146.810 104.075 147.545 ;
        RECT 104.345 147.375 104.515 147.545 ;
        RECT 105.260 147.495 105.975 147.665 ;
        RECT 106.170 147.545 106.490 147.835 ;
        RECT 106.665 147.545 107.005 148.515 ;
        RECT 107.175 147.545 107.345 148.685 ;
        RECT 107.615 147.885 107.865 148.685 ;
        RECT 108.510 147.715 108.840 148.515 ;
        RECT 109.140 147.885 109.470 148.685 ;
        RECT 109.640 147.715 109.970 148.515 ;
        RECT 107.535 147.545 109.970 147.715 ;
        RECT 110.345 147.595 112.015 148.685 ;
        RECT 112.185 147.925 112.700 148.335 ;
        RECT 112.935 147.925 113.105 148.685 ;
        RECT 113.275 148.345 115.305 148.515 ;
        RECT 104.245 147.045 104.515 147.375 ;
        RECT 104.685 147.045 105.090 147.375 ;
        RECT 105.260 147.045 105.970 147.495 ;
        RECT 104.345 146.875 104.515 147.045 ;
        RECT 103.905 146.465 104.175 146.810 ;
        RECT 104.345 146.705 105.955 146.875 ;
        RECT 106.140 146.805 106.490 147.375 ;
        RECT 106.665 146.985 106.840 147.545 ;
        RECT 107.535 147.295 107.705 147.545 ;
        RECT 107.010 147.125 107.705 147.295 ;
        RECT 107.880 147.125 108.300 147.325 ;
        RECT 108.470 147.125 108.800 147.325 ;
        RECT 108.970 147.125 109.300 147.325 ;
        RECT 106.665 146.935 106.895 146.985 ;
        RECT 104.365 146.135 104.745 146.535 ;
        RECT 104.915 146.355 105.085 146.705 ;
        RECT 105.255 146.135 105.585 146.535 ;
        RECT 105.785 146.355 105.955 146.705 ;
        RECT 106.155 146.135 106.485 146.635 ;
        RECT 106.665 146.305 107.005 146.935 ;
        RECT 107.175 146.135 107.425 146.935 ;
        RECT 107.615 146.785 108.840 146.955 ;
        RECT 107.615 146.305 107.945 146.785 ;
        RECT 108.115 146.135 108.340 146.595 ;
        RECT 108.510 146.305 108.840 146.785 ;
        RECT 109.470 146.915 109.640 147.545 ;
        RECT 109.825 147.125 110.175 147.375 ;
        RECT 110.345 147.075 111.095 147.595 ;
        RECT 109.470 146.305 109.970 146.915 ;
        RECT 111.265 146.905 112.015 147.425 ;
        RECT 112.185 147.115 112.525 147.925 ;
        RECT 113.275 147.680 113.445 148.345 ;
        RECT 113.840 148.005 114.965 148.175 ;
        RECT 112.695 147.490 113.445 147.680 ;
        RECT 113.615 147.665 114.625 147.835 ;
        RECT 112.185 146.945 113.415 147.115 ;
        RECT 110.345 146.135 112.015 146.905 ;
        RECT 112.460 146.340 112.705 146.945 ;
        RECT 112.925 146.135 113.435 146.670 ;
        RECT 113.615 146.305 113.805 147.665 ;
        RECT 113.975 147.325 114.250 147.465 ;
        RECT 113.975 147.155 114.255 147.325 ;
        RECT 113.975 146.305 114.250 147.155 ;
        RECT 114.455 146.865 114.625 147.665 ;
        RECT 114.795 146.875 114.965 148.005 ;
        RECT 115.135 147.375 115.305 148.345 ;
        RECT 115.475 147.545 115.645 148.685 ;
        RECT 115.815 147.545 116.150 148.515 ;
        RECT 115.135 147.045 115.330 147.375 ;
        RECT 115.555 147.045 115.810 147.375 ;
        RECT 115.555 146.875 115.725 147.045 ;
        RECT 115.980 146.875 116.150 147.545 ;
        RECT 116.700 147.705 116.955 148.375 ;
        RECT 117.135 147.885 117.420 148.685 ;
        RECT 117.600 147.965 117.930 148.475 ;
        RECT 116.700 146.985 116.880 147.705 ;
        RECT 117.600 147.375 117.850 147.965 ;
        RECT 118.200 147.815 118.370 148.425 ;
        RECT 118.540 147.995 118.870 148.685 ;
        RECT 119.100 148.135 119.340 148.425 ;
        RECT 119.540 148.305 119.960 148.685 ;
        RECT 120.140 148.215 120.770 148.465 ;
        RECT 121.240 148.305 121.570 148.685 ;
        RECT 120.140 148.135 120.310 148.215 ;
        RECT 121.740 148.135 121.910 148.425 ;
        RECT 122.090 148.305 122.470 148.685 ;
        RECT 122.710 148.300 123.540 148.470 ;
        RECT 119.100 147.965 120.310 148.135 ;
        RECT 117.050 147.045 117.850 147.375 ;
        RECT 114.795 146.705 115.725 146.875 ;
        RECT 114.795 146.670 114.970 146.705 ;
        RECT 114.440 146.305 114.970 146.670 ;
        RECT 115.395 146.135 115.725 146.535 ;
        RECT 115.895 146.305 116.150 146.875 ;
        RECT 116.615 146.845 116.880 146.985 ;
        RECT 116.615 146.815 116.955 146.845 ;
        RECT 116.700 146.315 116.955 146.815 ;
        RECT 117.135 146.135 117.420 146.595 ;
        RECT 117.600 146.395 117.850 147.045 ;
        RECT 118.050 147.795 118.370 147.815 ;
        RECT 118.050 147.625 119.970 147.795 ;
        RECT 118.050 146.730 118.240 147.625 ;
        RECT 120.140 147.455 120.310 147.965 ;
        RECT 120.480 147.705 121.000 148.015 ;
        RECT 118.410 147.285 120.310 147.455 ;
        RECT 118.410 147.225 118.740 147.285 ;
        RECT 118.890 147.055 119.220 147.115 ;
        RECT 118.560 146.785 119.220 147.055 ;
        RECT 118.050 146.400 118.370 146.730 ;
        RECT 118.550 146.135 119.210 146.615 ;
        RECT 119.410 146.525 119.580 147.285 ;
        RECT 120.480 147.115 120.660 147.525 ;
        RECT 119.750 146.945 120.080 147.065 ;
        RECT 120.830 146.945 121.000 147.705 ;
        RECT 119.750 146.775 121.000 146.945 ;
        RECT 121.170 147.885 122.540 148.135 ;
        RECT 121.170 147.115 121.360 147.885 ;
        RECT 122.290 147.625 122.540 147.885 ;
        RECT 121.530 147.455 121.780 147.615 ;
        RECT 122.710 147.455 122.880 148.300 ;
        RECT 123.775 148.015 123.945 148.515 ;
        RECT 124.115 148.185 124.445 148.685 ;
        RECT 123.050 147.625 123.550 148.005 ;
        RECT 123.775 147.845 124.470 148.015 ;
        RECT 121.530 147.285 122.880 147.455 ;
        RECT 122.460 147.245 122.880 147.285 ;
        RECT 121.170 146.775 121.590 147.115 ;
        RECT 121.880 146.785 122.290 147.115 ;
        RECT 119.410 146.355 120.260 146.525 ;
        RECT 120.820 146.135 121.140 146.595 ;
        RECT 121.340 146.345 121.590 146.775 ;
        RECT 121.880 146.135 122.290 146.575 ;
        RECT 122.460 146.515 122.630 147.245 ;
        RECT 122.800 146.695 123.150 147.065 ;
        RECT 123.330 146.755 123.550 147.625 ;
        RECT 123.720 147.055 124.130 147.675 ;
        RECT 124.300 146.875 124.470 147.845 ;
        RECT 123.775 146.685 124.470 146.875 ;
        RECT 122.460 146.315 123.475 146.515 ;
        RECT 123.775 146.355 123.945 146.685 ;
        RECT 124.115 146.135 124.445 146.515 ;
        RECT 124.660 146.395 124.885 148.515 ;
        RECT 125.055 148.185 125.385 148.685 ;
        RECT 125.555 148.015 125.725 148.515 ;
        RECT 125.060 147.845 125.725 148.015 ;
        RECT 125.060 146.855 125.290 147.845 ;
        RECT 125.460 147.025 125.810 147.675 ;
        RECT 126.445 147.595 127.655 148.685 ;
        RECT 126.445 147.055 126.965 147.595 ;
        RECT 127.135 146.885 127.655 147.425 ;
        RECT 125.060 146.685 125.725 146.855 ;
        RECT 125.055 146.135 125.385 146.515 ;
        RECT 125.555 146.395 125.725 146.685 ;
        RECT 126.445 146.135 127.655 146.885 ;
        RECT 14.580 145.965 127.740 146.135 ;
        RECT 14.665 145.215 15.875 145.965 ;
        RECT 14.665 144.675 15.185 145.215 ;
        RECT 16.045 145.195 19.555 145.965 ;
        RECT 15.355 144.505 15.875 145.045 ;
        RECT 14.665 143.415 15.875 144.505 ;
        RECT 16.045 144.505 17.735 145.025 ;
        RECT 17.905 144.675 19.555 145.195 ;
        RECT 19.765 145.145 19.995 145.965 ;
        RECT 20.165 145.165 20.495 145.795 ;
        RECT 19.745 144.725 20.075 144.975 ;
        RECT 20.245 144.565 20.495 145.165 ;
        RECT 20.665 145.145 20.875 145.965 ;
        RECT 21.145 145.145 21.375 145.965 ;
        RECT 21.545 145.165 21.875 145.795 ;
        RECT 21.125 144.725 21.455 144.975 ;
        RECT 21.625 144.565 21.875 145.165 ;
        RECT 22.045 145.145 22.255 145.965 ;
        RECT 22.860 145.625 23.115 145.785 ;
        RECT 22.775 145.455 23.115 145.625 ;
        RECT 23.295 145.505 23.580 145.965 ;
        RECT 22.860 145.255 23.115 145.455 ;
        RECT 16.045 143.415 19.555 144.505 ;
        RECT 19.765 143.415 19.995 144.555 ;
        RECT 20.165 143.585 20.495 144.565 ;
        RECT 20.665 143.415 20.875 144.555 ;
        RECT 21.145 143.415 21.375 144.555 ;
        RECT 21.545 143.585 21.875 144.565 ;
        RECT 22.045 143.415 22.255 144.555 ;
        RECT 22.860 144.395 23.040 145.255 ;
        RECT 23.760 145.055 24.010 145.705 ;
        RECT 23.210 144.725 24.010 145.055 ;
        RECT 22.860 143.725 23.115 144.395 ;
        RECT 23.295 143.415 23.580 144.215 ;
        RECT 23.760 144.135 24.010 144.725 ;
        RECT 24.210 145.370 24.530 145.700 ;
        RECT 24.710 145.485 25.370 145.965 ;
        RECT 25.570 145.575 26.420 145.745 ;
        RECT 24.210 144.475 24.400 145.370 ;
        RECT 24.720 145.045 25.380 145.315 ;
        RECT 25.050 144.985 25.380 145.045 ;
        RECT 24.570 144.815 24.900 144.875 ;
        RECT 25.570 144.815 25.740 145.575 ;
        RECT 26.980 145.505 27.300 145.965 ;
        RECT 27.500 145.325 27.750 145.755 ;
        RECT 28.040 145.525 28.450 145.965 ;
        RECT 28.620 145.585 29.635 145.785 ;
        RECT 25.910 145.155 27.160 145.325 ;
        RECT 25.910 145.035 26.240 145.155 ;
        RECT 24.570 144.645 26.470 144.815 ;
        RECT 24.210 144.305 26.130 144.475 ;
        RECT 24.210 144.285 24.530 144.305 ;
        RECT 23.760 143.625 24.090 144.135 ;
        RECT 24.360 143.675 24.530 144.285 ;
        RECT 26.300 144.135 26.470 144.645 ;
        RECT 26.640 144.575 26.820 144.985 ;
        RECT 26.990 144.395 27.160 145.155 ;
        RECT 24.700 143.415 25.030 144.105 ;
        RECT 25.260 143.965 26.470 144.135 ;
        RECT 26.640 144.085 27.160 144.395 ;
        RECT 27.330 144.985 27.750 145.325 ;
        RECT 28.040 144.985 28.450 145.315 ;
        RECT 27.330 144.215 27.520 144.985 ;
        RECT 28.620 144.855 28.790 145.585 ;
        RECT 29.935 145.415 30.105 145.745 ;
        RECT 30.275 145.585 30.605 145.965 ;
        RECT 28.960 145.035 29.310 145.405 ;
        RECT 28.620 144.815 29.040 144.855 ;
        RECT 27.690 144.645 29.040 144.815 ;
        RECT 27.690 144.485 27.940 144.645 ;
        RECT 28.450 144.215 28.700 144.475 ;
        RECT 27.330 143.965 28.700 144.215 ;
        RECT 25.260 143.675 25.500 143.965 ;
        RECT 26.300 143.885 26.470 143.965 ;
        RECT 25.700 143.415 26.120 143.795 ;
        RECT 26.300 143.635 26.930 143.885 ;
        RECT 27.400 143.415 27.730 143.795 ;
        RECT 27.900 143.675 28.070 143.965 ;
        RECT 28.870 143.800 29.040 144.645 ;
        RECT 29.490 144.475 29.710 145.345 ;
        RECT 29.935 145.225 30.630 145.415 ;
        RECT 29.210 144.095 29.710 144.475 ;
        RECT 29.880 144.425 30.290 145.045 ;
        RECT 30.460 144.255 30.630 145.225 ;
        RECT 29.935 144.085 30.630 144.255 ;
        RECT 28.250 143.415 28.630 143.795 ;
        RECT 28.870 143.630 29.700 143.800 ;
        RECT 29.935 143.585 30.105 144.085 ;
        RECT 30.275 143.415 30.605 143.915 ;
        RECT 30.820 143.585 31.045 145.705 ;
        RECT 31.215 145.585 31.545 145.965 ;
        RECT 31.715 145.415 31.885 145.705 ;
        RECT 31.220 145.245 31.885 145.415 ;
        RECT 31.220 144.255 31.450 145.245 ;
        RECT 32.145 145.215 33.355 145.965 ;
        RECT 31.620 144.425 31.970 145.075 ;
        RECT 32.145 144.505 32.665 145.045 ;
        RECT 32.835 144.675 33.355 145.215 ;
        RECT 33.525 145.195 37.035 145.965 ;
        RECT 37.205 145.240 37.495 145.965 ;
        RECT 38.125 145.195 40.715 145.965 ;
        RECT 33.525 144.505 35.215 145.025 ;
        RECT 35.385 144.675 37.035 145.195 ;
        RECT 31.220 144.085 31.885 144.255 ;
        RECT 31.215 143.415 31.545 143.915 ;
        RECT 31.715 143.585 31.885 144.085 ;
        RECT 32.145 143.415 33.355 144.505 ;
        RECT 33.525 143.415 37.035 144.505 ;
        RECT 37.205 143.415 37.495 144.580 ;
        RECT 38.125 144.505 39.335 145.025 ;
        RECT 39.505 144.675 40.715 145.195 ;
        RECT 40.925 145.145 41.155 145.965 ;
        RECT 41.325 145.165 41.655 145.795 ;
        RECT 40.905 144.725 41.235 144.975 ;
        RECT 41.405 144.565 41.655 145.165 ;
        RECT 41.825 145.145 42.035 145.965 ;
        RECT 42.640 145.255 42.895 145.785 ;
        RECT 43.075 145.505 43.360 145.965 ;
        RECT 42.640 144.605 42.820 145.255 ;
        RECT 43.540 145.055 43.790 145.705 ;
        RECT 42.990 144.725 43.790 145.055 ;
        RECT 38.125 143.415 40.715 144.505 ;
        RECT 40.925 143.415 41.155 144.555 ;
        RECT 41.325 143.585 41.655 144.565 ;
        RECT 41.825 143.415 42.035 144.555 ;
        RECT 42.555 144.435 42.820 144.605 ;
        RECT 42.640 144.395 42.820 144.435 ;
        RECT 42.640 143.725 42.895 144.395 ;
        RECT 43.075 143.415 43.360 144.215 ;
        RECT 43.540 144.135 43.790 144.725 ;
        RECT 43.990 145.370 44.310 145.700 ;
        RECT 44.490 145.485 45.150 145.965 ;
        RECT 45.350 145.575 46.200 145.745 ;
        RECT 43.990 144.475 44.180 145.370 ;
        RECT 44.500 145.045 45.160 145.315 ;
        RECT 44.830 144.985 45.160 145.045 ;
        RECT 44.350 144.815 44.680 144.875 ;
        RECT 45.350 144.815 45.520 145.575 ;
        RECT 46.760 145.505 47.080 145.965 ;
        RECT 47.280 145.325 47.530 145.755 ;
        RECT 47.820 145.525 48.230 145.965 ;
        RECT 48.400 145.585 49.415 145.785 ;
        RECT 45.690 145.155 46.940 145.325 ;
        RECT 45.690 145.035 46.020 145.155 ;
        RECT 44.350 144.645 46.250 144.815 ;
        RECT 43.990 144.305 45.910 144.475 ;
        RECT 43.990 144.285 44.310 144.305 ;
        RECT 43.540 143.625 43.870 144.135 ;
        RECT 44.140 143.675 44.310 144.285 ;
        RECT 46.080 144.135 46.250 144.645 ;
        RECT 46.420 144.575 46.600 144.985 ;
        RECT 46.770 144.395 46.940 145.155 ;
        RECT 44.480 143.415 44.810 144.105 ;
        RECT 45.040 143.965 46.250 144.135 ;
        RECT 46.420 144.085 46.940 144.395 ;
        RECT 47.110 144.985 47.530 145.325 ;
        RECT 47.820 144.985 48.230 145.315 ;
        RECT 47.110 144.215 47.300 144.985 ;
        RECT 48.400 144.855 48.570 145.585 ;
        RECT 49.715 145.415 49.885 145.745 ;
        RECT 50.055 145.585 50.385 145.965 ;
        RECT 48.740 145.035 49.090 145.405 ;
        RECT 48.400 144.815 48.820 144.855 ;
        RECT 47.470 144.645 48.820 144.815 ;
        RECT 47.470 144.485 47.720 144.645 ;
        RECT 48.230 144.215 48.480 144.475 ;
        RECT 47.110 143.965 48.480 144.215 ;
        RECT 45.040 143.675 45.280 143.965 ;
        RECT 46.080 143.885 46.250 143.965 ;
        RECT 45.480 143.415 45.900 143.795 ;
        RECT 46.080 143.635 46.710 143.885 ;
        RECT 47.180 143.415 47.510 143.795 ;
        RECT 47.680 143.675 47.850 143.965 ;
        RECT 48.650 143.800 48.820 144.645 ;
        RECT 49.270 144.475 49.490 145.345 ;
        RECT 49.715 145.225 50.410 145.415 ;
        RECT 48.990 144.095 49.490 144.475 ;
        RECT 49.660 144.425 50.070 145.045 ;
        RECT 50.240 144.255 50.410 145.225 ;
        RECT 49.715 144.085 50.410 144.255 ;
        RECT 48.030 143.415 48.410 143.795 ;
        RECT 48.650 143.630 49.480 143.800 ;
        RECT 49.715 143.585 49.885 144.085 ;
        RECT 50.055 143.415 50.385 143.915 ;
        RECT 50.600 143.585 50.825 145.705 ;
        RECT 50.995 145.585 51.325 145.965 ;
        RECT 51.495 145.415 51.665 145.705 ;
        RECT 51.000 145.245 51.665 145.415 ;
        RECT 51.000 144.255 51.230 145.245 ;
        RECT 51.930 145.225 52.185 145.795 ;
        RECT 52.355 145.565 52.685 145.965 ;
        RECT 53.110 145.430 53.640 145.795 ;
        RECT 53.830 145.625 54.105 145.795 ;
        RECT 53.825 145.455 54.105 145.625 ;
        RECT 53.110 145.395 53.285 145.430 ;
        RECT 52.355 145.225 53.285 145.395 ;
        RECT 51.400 144.425 51.750 145.075 ;
        RECT 51.930 144.555 52.100 145.225 ;
        RECT 52.355 145.055 52.525 145.225 ;
        RECT 52.270 144.725 52.525 145.055 ;
        RECT 52.750 144.725 52.945 145.055 ;
        RECT 51.000 144.085 51.665 144.255 ;
        RECT 50.995 143.415 51.325 143.915 ;
        RECT 51.495 143.585 51.665 144.085 ;
        RECT 51.930 143.585 52.265 144.555 ;
        RECT 52.435 143.415 52.605 144.555 ;
        RECT 52.775 143.755 52.945 144.725 ;
        RECT 53.115 144.095 53.285 145.225 ;
        RECT 53.455 144.435 53.625 145.235 ;
        RECT 53.830 144.635 54.105 145.455 ;
        RECT 54.275 144.435 54.465 145.795 ;
        RECT 54.645 145.430 55.155 145.965 ;
        RECT 55.375 145.155 55.620 145.760 ;
        RECT 56.525 145.195 58.195 145.965 ;
        RECT 54.665 144.985 55.895 145.155 ;
        RECT 53.455 144.265 54.465 144.435 ;
        RECT 54.635 144.420 55.385 144.610 ;
        RECT 53.115 143.925 54.240 144.095 ;
        RECT 54.635 143.755 54.805 144.420 ;
        RECT 55.555 144.175 55.895 144.985 ;
        RECT 52.775 143.585 54.805 143.755 ;
        RECT 54.975 143.415 55.145 144.175 ;
        RECT 55.380 143.765 55.895 144.175 ;
        RECT 56.525 144.505 57.275 145.025 ;
        RECT 57.445 144.675 58.195 145.195 ;
        RECT 58.405 145.145 58.635 145.965 ;
        RECT 58.805 145.165 59.135 145.795 ;
        RECT 58.385 144.725 58.715 144.975 ;
        RECT 58.885 144.565 59.135 145.165 ;
        RECT 59.305 145.145 59.515 145.965 ;
        RECT 60.205 145.195 62.795 145.965 ;
        RECT 62.965 145.240 63.255 145.965 ;
        RECT 56.525 143.415 58.195 144.505 ;
        RECT 58.405 143.415 58.635 144.555 ;
        RECT 58.805 143.585 59.135 144.565 ;
        RECT 59.305 143.415 59.515 144.555 ;
        RECT 60.205 144.505 61.415 145.025 ;
        RECT 61.585 144.675 62.795 145.195 ;
        RECT 64.160 145.155 64.405 145.760 ;
        RECT 64.625 145.430 65.135 145.965 ;
        RECT 63.885 144.985 65.115 145.155 ;
        RECT 60.205 143.415 62.795 144.505 ;
        RECT 62.965 143.415 63.255 144.580 ;
        RECT 63.885 144.175 64.225 144.985 ;
        RECT 64.395 144.420 65.145 144.610 ;
        RECT 63.885 143.765 64.400 144.175 ;
        RECT 64.635 143.415 64.805 144.175 ;
        RECT 64.975 143.755 65.145 144.420 ;
        RECT 65.315 144.435 65.505 145.795 ;
        RECT 65.675 144.945 65.950 145.795 ;
        RECT 66.140 145.430 66.670 145.795 ;
        RECT 67.095 145.565 67.425 145.965 ;
        RECT 66.495 145.395 66.670 145.430 ;
        RECT 65.675 144.775 65.955 144.945 ;
        RECT 65.675 144.635 65.950 144.775 ;
        RECT 66.155 144.435 66.325 145.235 ;
        RECT 65.315 144.265 66.325 144.435 ;
        RECT 66.495 145.225 67.425 145.395 ;
        RECT 67.595 145.225 67.850 145.795 ;
        RECT 68.490 145.420 73.835 145.965 ;
        RECT 74.010 145.420 79.355 145.965 ;
        RECT 79.535 145.465 79.865 145.965 ;
        RECT 66.495 144.095 66.665 145.225 ;
        RECT 67.255 145.055 67.425 145.225 ;
        RECT 65.540 143.925 66.665 144.095 ;
        RECT 66.835 144.725 67.030 145.055 ;
        RECT 67.255 144.725 67.510 145.055 ;
        RECT 66.835 143.755 67.005 144.725 ;
        RECT 67.680 144.555 67.850 145.225 ;
        RECT 64.975 143.585 67.005 143.755 ;
        RECT 67.175 143.415 67.345 144.555 ;
        RECT 67.515 143.585 67.850 144.555 ;
        RECT 70.080 143.850 70.430 145.100 ;
        RECT 71.910 144.590 72.250 145.420 ;
        RECT 75.600 143.850 75.950 145.100 ;
        RECT 77.430 144.590 77.770 145.420 ;
        RECT 80.065 145.395 80.235 145.745 ;
        RECT 80.435 145.565 80.765 145.965 ;
        RECT 80.935 145.395 81.105 145.745 ;
        RECT 81.275 145.565 81.655 145.965 ;
        RECT 79.530 144.725 79.880 145.295 ;
        RECT 80.065 145.225 81.675 145.395 ;
        RECT 81.845 145.290 82.115 145.635 ;
        RECT 81.505 145.055 81.675 145.225 ;
        RECT 79.530 144.265 79.850 144.555 ;
        RECT 80.050 144.435 80.760 145.055 ;
        RECT 80.930 144.725 81.335 145.055 ;
        RECT 81.505 144.725 81.775 145.055 ;
        RECT 81.505 144.555 81.675 144.725 ;
        RECT 81.945 144.555 82.115 145.290 ;
        RECT 82.745 145.195 84.415 145.965 ;
        RECT 80.950 144.385 81.675 144.555 ;
        RECT 80.950 144.265 81.120 144.385 ;
        RECT 79.530 144.095 81.120 144.265 ;
        RECT 68.490 143.415 73.835 143.850 ;
        RECT 74.010 143.415 79.355 143.850 ;
        RECT 79.530 143.635 81.185 143.925 ;
        RECT 81.355 143.415 81.635 144.215 ;
        RECT 81.845 143.585 82.115 144.555 ;
        RECT 82.745 144.505 83.495 145.025 ;
        RECT 83.665 144.675 84.415 145.195 ;
        RECT 84.860 145.155 85.105 145.760 ;
        RECT 85.325 145.430 85.835 145.965 ;
        RECT 84.585 144.985 85.815 145.155 ;
        RECT 82.745 143.415 84.415 144.505 ;
        RECT 84.585 144.175 84.925 144.985 ;
        RECT 85.095 144.420 85.845 144.610 ;
        RECT 84.585 143.765 85.100 144.175 ;
        RECT 85.335 143.415 85.505 144.175 ;
        RECT 85.675 143.755 85.845 144.420 ;
        RECT 86.015 144.435 86.205 145.795 ;
        RECT 86.375 144.945 86.650 145.795 ;
        RECT 86.840 145.430 87.370 145.795 ;
        RECT 87.795 145.565 88.125 145.965 ;
        RECT 87.195 145.395 87.370 145.430 ;
        RECT 86.375 144.775 86.655 144.945 ;
        RECT 86.375 144.635 86.650 144.775 ;
        RECT 86.855 144.435 87.025 145.235 ;
        RECT 86.015 144.265 87.025 144.435 ;
        RECT 87.195 145.225 88.125 145.395 ;
        RECT 88.295 145.225 88.550 145.795 ;
        RECT 88.725 145.240 89.015 145.965 ;
        RECT 90.195 145.415 90.365 145.795 ;
        RECT 90.545 145.585 90.875 145.965 ;
        RECT 90.195 145.245 90.860 145.415 ;
        RECT 91.055 145.290 91.315 145.795 ;
        RECT 87.195 144.095 87.365 145.225 ;
        RECT 87.955 145.055 88.125 145.225 ;
        RECT 86.240 143.925 87.365 144.095 ;
        RECT 87.535 144.725 87.730 145.055 ;
        RECT 87.955 144.725 88.210 145.055 ;
        RECT 87.535 143.755 87.705 144.725 ;
        RECT 88.380 144.555 88.550 145.225 ;
        RECT 90.125 144.695 90.455 145.065 ;
        RECT 90.690 144.990 90.860 145.245 ;
        RECT 90.690 144.660 90.975 144.990 ;
        RECT 85.675 143.585 87.705 143.755 ;
        RECT 87.875 143.415 88.045 144.555 ;
        RECT 88.215 143.585 88.550 144.555 ;
        RECT 88.725 143.415 89.015 144.580 ;
        RECT 90.690 144.515 90.860 144.660 ;
        RECT 90.195 144.345 90.860 144.515 ;
        RECT 91.145 144.490 91.315 145.290 ;
        RECT 91.945 145.195 93.615 145.965 ;
        RECT 90.195 143.585 90.365 144.345 ;
        RECT 90.545 143.415 90.875 144.175 ;
        RECT 91.045 143.585 91.315 144.490 ;
        RECT 91.945 144.505 92.695 145.025 ;
        RECT 92.865 144.675 93.615 145.195 ;
        RECT 93.900 145.335 94.185 145.795 ;
        RECT 94.355 145.505 94.625 145.965 ;
        RECT 93.900 145.165 94.855 145.335 ;
        RECT 91.945 143.415 93.615 144.505 ;
        RECT 93.785 144.435 94.475 144.995 ;
        RECT 94.645 144.265 94.855 145.165 ;
        RECT 93.900 144.045 94.855 144.265 ;
        RECT 95.025 144.995 95.425 145.795 ;
        RECT 95.615 145.335 95.895 145.795 ;
        RECT 96.415 145.505 96.740 145.965 ;
        RECT 95.615 145.165 96.740 145.335 ;
        RECT 96.910 145.225 97.295 145.795 ;
        RECT 96.290 145.055 96.740 145.165 ;
        RECT 95.025 144.435 96.120 144.995 ;
        RECT 96.290 144.725 96.845 145.055 ;
        RECT 93.900 143.585 94.185 144.045 ;
        RECT 94.355 143.415 94.625 143.875 ;
        RECT 95.025 143.585 95.425 144.435 ;
        RECT 96.290 144.265 96.740 144.725 ;
        RECT 97.015 144.555 97.295 145.225 ;
        RECT 97.925 145.195 101.435 145.965 ;
        RECT 101.610 145.420 106.955 145.965 ;
        RECT 107.135 145.465 107.465 145.965 ;
        RECT 95.615 144.045 96.740 144.265 ;
        RECT 95.615 143.585 95.895 144.045 ;
        RECT 96.415 143.415 96.740 143.875 ;
        RECT 96.910 143.585 97.295 144.555 ;
        RECT 97.925 144.505 99.615 145.025 ;
        RECT 99.785 144.675 101.435 145.195 ;
        RECT 97.925 143.415 101.435 144.505 ;
        RECT 103.200 143.850 103.550 145.100 ;
        RECT 105.030 144.590 105.370 145.420 ;
        RECT 107.665 145.395 107.835 145.745 ;
        RECT 108.035 145.565 108.365 145.965 ;
        RECT 108.535 145.395 108.705 145.745 ;
        RECT 108.875 145.565 109.255 145.965 ;
        RECT 107.130 144.725 107.480 145.295 ;
        RECT 107.665 145.225 109.275 145.395 ;
        RECT 109.445 145.290 109.715 145.635 ;
        RECT 109.105 145.055 109.275 145.225 ;
        RECT 107.130 144.265 107.450 144.555 ;
        RECT 107.650 144.435 108.360 145.055 ;
        RECT 108.530 144.725 108.935 145.055 ;
        RECT 109.105 144.725 109.375 145.055 ;
        RECT 109.105 144.555 109.275 144.725 ;
        RECT 109.545 144.555 109.715 145.290 ;
        RECT 108.550 144.385 109.275 144.555 ;
        RECT 108.550 144.265 108.720 144.385 ;
        RECT 107.130 144.095 108.720 144.265 ;
        RECT 101.610 143.415 106.955 143.850 ;
        RECT 107.130 143.635 108.785 143.925 ;
        RECT 108.955 143.415 109.235 144.215 ;
        RECT 109.445 143.585 109.715 144.555 ;
        RECT 109.885 145.165 110.225 145.795 ;
        RECT 110.395 145.165 110.645 145.965 ;
        RECT 110.835 145.315 111.165 145.795 ;
        RECT 111.335 145.505 111.560 145.965 ;
        RECT 111.730 145.315 112.060 145.795 ;
        RECT 109.885 145.115 110.115 145.165 ;
        RECT 110.835 145.145 112.060 145.315 ;
        RECT 112.690 145.185 113.190 145.795 ;
        RECT 114.485 145.240 114.775 145.965 ;
        RECT 109.885 144.555 110.060 145.115 ;
        RECT 110.230 144.805 110.925 144.975 ;
        RECT 110.755 144.555 110.925 144.805 ;
        RECT 111.100 144.775 111.520 144.975 ;
        RECT 111.690 144.775 112.020 144.975 ;
        RECT 112.190 144.775 112.520 144.975 ;
        RECT 112.690 144.555 112.860 145.185 ;
        RECT 115.680 145.155 115.925 145.760 ;
        RECT 116.145 145.430 116.655 145.965 ;
        RECT 115.405 144.985 116.635 145.155 ;
        RECT 113.045 144.725 113.395 144.975 ;
        RECT 109.885 143.585 110.225 144.555 ;
        RECT 110.395 143.415 110.565 144.555 ;
        RECT 110.755 144.385 113.190 144.555 ;
        RECT 110.835 143.415 111.085 144.215 ;
        RECT 111.730 143.585 112.060 144.385 ;
        RECT 112.360 143.415 112.690 144.215 ;
        RECT 112.860 143.585 113.190 144.385 ;
        RECT 114.485 143.415 114.775 144.580 ;
        RECT 115.405 144.175 115.745 144.985 ;
        RECT 115.915 144.420 116.665 144.610 ;
        RECT 115.405 143.765 115.920 144.175 ;
        RECT 116.155 143.415 116.325 144.175 ;
        RECT 116.495 143.755 116.665 144.420 ;
        RECT 116.835 144.435 117.025 145.795 ;
        RECT 117.195 145.625 117.470 145.795 ;
        RECT 117.195 145.455 117.475 145.625 ;
        RECT 117.195 144.635 117.470 145.455 ;
        RECT 117.660 145.430 118.190 145.795 ;
        RECT 118.615 145.565 118.945 145.965 ;
        RECT 118.015 145.395 118.190 145.430 ;
        RECT 117.675 144.435 117.845 145.235 ;
        RECT 116.835 144.265 117.845 144.435 ;
        RECT 118.015 145.225 118.945 145.395 ;
        RECT 119.115 145.225 119.370 145.795 ;
        RECT 118.015 144.095 118.185 145.225 ;
        RECT 118.775 145.055 118.945 145.225 ;
        RECT 117.060 143.925 118.185 144.095 ;
        RECT 118.355 144.725 118.550 145.055 ;
        RECT 118.775 144.725 119.030 145.055 ;
        RECT 118.355 143.755 118.525 144.725 ;
        RECT 119.200 144.555 119.370 145.225 ;
        RECT 119.585 145.145 119.815 145.965 ;
        RECT 119.985 145.165 120.315 145.795 ;
        RECT 119.565 144.725 119.895 144.975 ;
        RECT 120.065 144.565 120.315 145.165 ;
        RECT 120.485 145.145 120.695 145.965 ;
        RECT 121.475 145.415 121.645 145.795 ;
        RECT 121.825 145.585 122.155 145.965 ;
        RECT 121.475 145.245 122.140 145.415 ;
        RECT 122.335 145.290 122.595 145.795 ;
        RECT 121.405 144.695 121.735 145.065 ;
        RECT 121.970 144.990 122.140 145.245 ;
        RECT 116.495 143.585 118.525 143.755 ;
        RECT 118.695 143.415 118.865 144.555 ;
        RECT 119.035 143.585 119.370 144.555 ;
        RECT 119.585 143.415 119.815 144.555 ;
        RECT 119.985 143.585 120.315 144.565 ;
        RECT 121.970 144.660 122.255 144.990 ;
        RECT 120.485 143.415 120.695 144.555 ;
        RECT 121.970 144.515 122.140 144.660 ;
        RECT 121.475 144.345 122.140 144.515 ;
        RECT 122.425 144.490 122.595 145.290 ;
        RECT 122.765 145.195 126.275 145.965 ;
        RECT 126.445 145.215 127.655 145.965 ;
        RECT 121.475 143.585 121.645 144.345 ;
        RECT 121.825 143.415 122.155 144.175 ;
        RECT 122.325 143.585 122.595 144.490 ;
        RECT 122.765 144.505 124.455 145.025 ;
        RECT 124.625 144.675 126.275 145.195 ;
        RECT 126.445 144.505 126.965 145.045 ;
        RECT 127.135 144.675 127.655 145.215 ;
        RECT 122.765 143.415 126.275 144.505 ;
        RECT 126.445 143.415 127.655 144.505 ;
        RECT 14.580 143.245 127.740 143.415 ;
        RECT 14.665 142.155 15.875 143.245 ;
        RECT 14.665 141.445 15.185 141.985 ;
        RECT 15.355 141.615 15.875 142.155 ;
        RECT 16.045 142.155 18.635 143.245 ;
        RECT 18.810 142.810 24.155 143.245 ;
        RECT 16.045 141.635 17.255 142.155 ;
        RECT 17.425 141.465 18.635 141.985 ;
        RECT 20.400 141.560 20.750 142.810 ;
        RECT 24.325 142.080 24.615 143.245 ;
        RECT 25.245 142.155 28.755 143.245 ;
        RECT 28.930 142.810 34.275 143.245 ;
        RECT 14.665 140.695 15.875 141.445 ;
        RECT 16.045 140.695 18.635 141.465 ;
        RECT 22.230 141.240 22.570 142.070 ;
        RECT 25.245 141.635 26.935 142.155 ;
        RECT 27.105 141.465 28.755 141.985 ;
        RECT 30.520 141.560 30.870 142.810 ;
        RECT 34.445 142.105 34.715 143.075 ;
        RECT 34.925 142.445 35.205 143.245 ;
        RECT 35.375 142.735 37.030 143.025 ;
        RECT 35.440 142.395 37.030 142.565 ;
        RECT 35.440 142.275 35.610 142.395 ;
        RECT 34.885 142.105 35.610 142.275 ;
        RECT 18.810 140.695 24.155 141.240 ;
        RECT 24.325 140.695 24.615 141.420 ;
        RECT 25.245 140.695 28.755 141.465 ;
        RECT 32.350 141.240 32.690 142.070 ;
        RECT 34.445 141.370 34.615 142.105 ;
        RECT 34.885 141.935 35.055 142.105 ;
        RECT 34.785 141.605 35.055 141.935 ;
        RECT 35.225 141.605 35.630 141.935 ;
        RECT 35.800 141.605 36.510 142.225 ;
        RECT 36.710 142.105 37.030 142.395 ;
        RECT 38.125 142.155 41.635 143.245 ;
        RECT 41.810 142.810 47.155 143.245 ;
        RECT 34.885 141.435 35.055 141.605 ;
        RECT 28.930 140.695 34.275 141.240 ;
        RECT 34.445 141.025 34.715 141.370 ;
        RECT 34.885 141.265 36.495 141.435 ;
        RECT 36.680 141.365 37.030 141.935 ;
        RECT 38.125 141.635 39.815 142.155 ;
        RECT 39.985 141.465 41.635 141.985 ;
        RECT 43.400 141.560 43.750 142.810 ;
        RECT 47.325 142.105 47.595 143.075 ;
        RECT 47.805 142.445 48.085 143.245 ;
        RECT 48.255 142.735 49.910 143.025 ;
        RECT 48.320 142.395 49.910 142.565 ;
        RECT 48.320 142.275 48.490 142.395 ;
        RECT 47.765 142.105 48.490 142.275 ;
        RECT 34.905 140.695 35.285 141.095 ;
        RECT 35.455 140.915 35.625 141.265 ;
        RECT 35.795 140.695 36.125 141.095 ;
        RECT 36.325 140.915 36.495 141.265 ;
        RECT 36.695 140.695 37.025 141.195 ;
        RECT 38.125 140.695 41.635 141.465 ;
        RECT 45.230 141.240 45.570 142.070 ;
        RECT 47.325 141.370 47.495 142.105 ;
        RECT 47.765 141.935 47.935 142.105 ;
        RECT 47.665 141.605 47.935 141.935 ;
        RECT 48.105 141.605 48.510 141.935 ;
        RECT 48.680 141.605 49.390 142.225 ;
        RECT 49.590 142.105 49.910 142.395 ;
        RECT 50.085 142.080 50.375 143.245 ;
        RECT 50.545 142.155 52.215 143.245 ;
        RECT 47.765 141.435 47.935 141.605 ;
        RECT 41.810 140.695 47.155 141.240 ;
        RECT 47.325 141.025 47.595 141.370 ;
        RECT 47.765 141.265 49.375 141.435 ;
        RECT 49.560 141.365 49.910 141.935 ;
        RECT 50.545 141.635 51.295 142.155 ;
        RECT 52.385 142.105 52.725 143.075 ;
        RECT 52.895 142.105 53.065 143.245 ;
        RECT 53.335 142.445 53.585 143.245 ;
        RECT 54.230 142.275 54.560 143.075 ;
        RECT 54.860 142.445 55.190 143.245 ;
        RECT 55.360 142.275 55.690 143.075 ;
        RECT 56.180 142.615 56.465 143.075 ;
        RECT 56.635 142.785 56.905 143.245 ;
        RECT 56.180 142.395 57.135 142.615 ;
        RECT 53.255 142.105 55.690 142.275 ;
        RECT 51.465 141.465 52.215 141.985 ;
        RECT 47.785 140.695 48.165 141.095 ;
        RECT 48.335 140.915 48.505 141.265 ;
        RECT 48.675 140.695 49.005 141.095 ;
        RECT 49.205 140.915 49.375 141.265 ;
        RECT 49.575 140.695 49.905 141.195 ;
        RECT 50.085 140.695 50.375 141.420 ;
        RECT 50.545 140.695 52.215 141.465 ;
        RECT 52.385 141.545 52.560 142.105 ;
        RECT 53.255 141.855 53.425 142.105 ;
        RECT 52.730 141.685 53.425 141.855 ;
        RECT 53.600 141.685 54.020 141.885 ;
        RECT 54.190 141.685 54.520 141.885 ;
        RECT 54.690 141.685 55.020 141.885 ;
        RECT 52.385 141.495 52.615 141.545 ;
        RECT 52.385 140.865 52.725 141.495 ;
        RECT 52.895 140.695 53.145 141.495 ;
        RECT 53.335 141.345 54.560 141.515 ;
        RECT 53.335 140.865 53.665 141.345 ;
        RECT 53.835 140.695 54.060 141.155 ;
        RECT 54.230 140.865 54.560 141.345 ;
        RECT 55.190 141.475 55.360 142.105 ;
        RECT 55.545 141.685 55.895 141.935 ;
        RECT 56.065 141.665 56.755 142.225 ;
        RECT 56.925 141.495 57.135 142.395 ;
        RECT 55.190 140.865 55.690 141.475 ;
        RECT 56.180 141.325 57.135 141.495 ;
        RECT 57.305 142.225 57.705 143.075 ;
        RECT 57.895 142.615 58.175 143.075 ;
        RECT 58.695 142.785 59.020 143.245 ;
        RECT 57.895 142.395 59.020 142.615 ;
        RECT 57.305 141.665 58.400 142.225 ;
        RECT 58.570 141.935 59.020 142.395 ;
        RECT 59.190 142.105 59.575 143.075 ;
        RECT 56.180 140.865 56.465 141.325 ;
        RECT 56.635 140.695 56.905 141.155 ;
        RECT 57.305 140.865 57.705 141.665 ;
        RECT 58.570 141.605 59.125 141.935 ;
        RECT 58.570 141.495 59.020 141.605 ;
        RECT 57.895 141.325 59.020 141.495 ;
        RECT 59.295 141.435 59.575 142.105 ;
        RECT 57.895 140.865 58.175 141.325 ;
        RECT 58.695 140.695 59.020 141.155 ;
        RECT 59.190 140.865 59.575 141.435 ;
        RECT 59.750 142.055 60.005 142.935 ;
        RECT 60.175 142.105 60.480 143.245 ;
        RECT 60.820 142.865 61.150 143.245 ;
        RECT 61.330 142.695 61.500 142.985 ;
        RECT 61.670 142.785 61.920 143.245 ;
        RECT 60.700 142.525 61.500 142.695 ;
        RECT 62.090 142.735 62.960 143.075 ;
        RECT 59.750 141.405 59.960 142.055 ;
        RECT 60.700 141.935 60.870 142.525 ;
        RECT 62.090 142.355 62.260 142.735 ;
        RECT 63.195 142.615 63.365 143.075 ;
        RECT 63.535 142.785 63.905 143.245 ;
        RECT 64.200 142.645 64.370 142.985 ;
        RECT 64.540 142.815 64.870 143.245 ;
        RECT 65.105 142.645 65.275 142.985 ;
        RECT 61.040 142.185 62.260 142.355 ;
        RECT 62.430 142.275 62.890 142.565 ;
        RECT 63.195 142.445 63.755 142.615 ;
        RECT 64.200 142.475 65.275 142.645 ;
        RECT 65.445 142.745 66.125 143.075 ;
        RECT 66.340 142.745 66.590 143.075 ;
        RECT 66.760 142.785 67.010 143.245 ;
        RECT 63.585 142.305 63.755 142.445 ;
        RECT 62.430 142.265 63.395 142.275 ;
        RECT 62.090 142.095 62.260 142.185 ;
        RECT 62.720 142.105 63.395 142.265 ;
        RECT 60.130 141.905 60.870 141.935 ;
        RECT 60.130 141.605 61.045 141.905 ;
        RECT 60.720 141.430 61.045 141.605 ;
        RECT 59.750 140.875 60.005 141.405 ;
        RECT 60.175 140.695 60.480 141.155 ;
        RECT 60.725 141.075 61.045 141.430 ;
        RECT 61.215 141.645 61.755 142.015 ;
        RECT 62.090 141.925 62.495 142.095 ;
        RECT 61.215 141.245 61.455 141.645 ;
        RECT 61.935 141.475 62.155 141.755 ;
        RECT 61.625 141.305 62.155 141.475 ;
        RECT 61.625 141.075 61.795 141.305 ;
        RECT 62.325 141.145 62.495 141.925 ;
        RECT 62.665 141.315 63.015 141.935 ;
        RECT 63.185 141.315 63.395 142.105 ;
        RECT 63.585 142.135 65.085 142.305 ;
        RECT 63.585 141.445 63.755 142.135 ;
        RECT 65.445 141.965 65.615 142.745 ;
        RECT 66.420 142.615 66.590 142.745 ;
        RECT 63.925 141.795 65.615 141.965 ;
        RECT 65.785 142.185 66.250 142.575 ;
        RECT 66.420 142.445 66.815 142.615 ;
        RECT 63.925 141.615 64.095 141.795 ;
        RECT 60.725 140.905 61.795 141.075 ;
        RECT 61.965 140.695 62.155 141.135 ;
        RECT 62.325 140.865 63.275 141.145 ;
        RECT 63.585 141.055 63.845 141.445 ;
        RECT 64.265 141.375 65.055 141.625 ;
        RECT 63.495 140.885 63.845 141.055 ;
        RECT 64.055 140.695 64.385 141.155 ;
        RECT 65.260 141.085 65.430 141.795 ;
        RECT 65.785 141.595 65.955 142.185 ;
        RECT 65.600 141.375 65.955 141.595 ;
        RECT 66.125 141.375 66.475 141.995 ;
        RECT 66.645 141.085 66.815 142.445 ;
        RECT 67.180 142.275 67.505 143.060 ;
        RECT 66.985 141.225 67.445 142.275 ;
        RECT 65.260 140.915 66.115 141.085 ;
        RECT 66.320 140.915 66.815 141.085 ;
        RECT 66.985 140.695 67.315 141.055 ;
        RECT 67.675 140.955 67.845 143.075 ;
        RECT 68.015 142.745 68.345 143.245 ;
        RECT 68.515 142.575 68.770 143.075 ;
        RECT 68.020 142.405 68.770 142.575 ;
        RECT 68.020 141.415 68.250 142.405 ;
        RECT 68.420 141.585 68.770 142.235 ;
        RECT 68.945 142.170 69.215 143.075 ;
        RECT 69.385 142.485 69.715 143.245 ;
        RECT 69.895 142.315 70.065 143.075 ;
        RECT 68.020 141.245 68.770 141.415 ;
        RECT 68.015 140.695 68.345 141.075 ;
        RECT 68.515 140.955 68.770 141.245 ;
        RECT 68.945 141.370 69.115 142.170 ;
        RECT 69.400 142.145 70.065 142.315 ;
        RECT 70.325 142.155 71.535 143.245 ;
        RECT 69.400 142.000 69.570 142.145 ;
        RECT 69.285 141.670 69.570 142.000 ;
        RECT 69.400 141.415 69.570 141.670 ;
        RECT 69.805 141.595 70.135 141.965 ;
        RECT 70.325 141.615 70.845 142.155 ;
        RECT 71.765 142.105 71.975 143.245 ;
        RECT 72.145 142.095 72.475 143.075 ;
        RECT 72.645 142.105 72.875 143.245 ;
        RECT 73.085 142.155 75.675 143.245 ;
        RECT 71.015 141.445 71.535 141.985 ;
        RECT 68.945 140.865 69.205 141.370 ;
        RECT 69.400 141.245 70.065 141.415 ;
        RECT 69.385 140.695 69.715 141.075 ;
        RECT 69.895 140.865 70.065 141.245 ;
        RECT 70.325 140.695 71.535 141.445 ;
        RECT 71.765 140.695 71.975 141.515 ;
        RECT 72.145 141.495 72.395 142.095 ;
        RECT 72.565 141.685 72.895 141.935 ;
        RECT 73.085 141.635 74.295 142.155 ;
        RECT 75.845 142.080 76.135 143.245 ;
        RECT 76.765 142.155 79.355 143.245 ;
        RECT 79.530 142.810 84.875 143.245 ;
        RECT 85.050 142.810 90.395 143.245 ;
        RECT 90.570 142.810 95.915 143.245 ;
        RECT 96.090 142.810 101.435 143.245 ;
        RECT 72.145 140.865 72.475 141.495 ;
        RECT 72.645 140.695 72.875 141.515 ;
        RECT 74.465 141.465 75.675 141.985 ;
        RECT 76.765 141.635 77.975 142.155 ;
        RECT 78.145 141.465 79.355 141.985 ;
        RECT 81.120 141.560 81.470 142.810 ;
        RECT 73.085 140.695 75.675 141.465 ;
        RECT 75.845 140.695 76.135 141.420 ;
        RECT 76.765 140.695 79.355 141.465 ;
        RECT 82.950 141.240 83.290 142.070 ;
        RECT 86.640 141.560 86.990 142.810 ;
        RECT 88.470 141.240 88.810 142.070 ;
        RECT 92.160 141.560 92.510 142.810 ;
        RECT 93.990 141.240 94.330 142.070 ;
        RECT 97.680 141.560 98.030 142.810 ;
        RECT 101.605 142.080 101.895 143.245 ;
        RECT 102.065 142.155 104.655 143.245 ;
        RECT 104.830 142.810 110.175 143.245 ;
        RECT 110.350 142.810 115.695 143.245 ;
        RECT 99.510 141.240 99.850 142.070 ;
        RECT 102.065 141.635 103.275 142.155 ;
        RECT 103.445 141.465 104.655 141.985 ;
        RECT 106.420 141.560 106.770 142.810 ;
        RECT 79.530 140.695 84.875 141.240 ;
        RECT 85.050 140.695 90.395 141.240 ;
        RECT 90.570 140.695 95.915 141.240 ;
        RECT 96.090 140.695 101.435 141.240 ;
        RECT 101.605 140.695 101.895 141.420 ;
        RECT 102.065 140.695 104.655 141.465 ;
        RECT 108.250 141.240 108.590 142.070 ;
        RECT 111.940 141.560 112.290 142.810 ;
        RECT 115.865 142.485 116.380 142.895 ;
        RECT 116.615 142.485 116.785 143.245 ;
        RECT 116.955 142.905 118.985 143.075 ;
        RECT 113.770 141.240 114.110 142.070 ;
        RECT 115.865 141.675 116.205 142.485 ;
        RECT 116.955 142.240 117.125 142.905 ;
        RECT 117.520 142.565 118.645 142.735 ;
        RECT 116.375 142.050 117.125 142.240 ;
        RECT 117.295 142.225 118.305 142.395 ;
        RECT 115.865 141.505 117.095 141.675 ;
        RECT 104.830 140.695 110.175 141.240 ;
        RECT 110.350 140.695 115.695 141.240 ;
        RECT 116.140 140.900 116.385 141.505 ;
        RECT 116.605 140.695 117.115 141.230 ;
        RECT 117.295 140.865 117.485 142.225 ;
        RECT 117.655 141.885 117.930 142.025 ;
        RECT 117.655 141.715 117.935 141.885 ;
        RECT 117.655 140.865 117.930 141.715 ;
        RECT 118.135 141.425 118.305 142.225 ;
        RECT 118.475 141.435 118.645 142.565 ;
        RECT 118.815 141.935 118.985 142.905 ;
        RECT 119.155 142.105 119.325 143.245 ;
        RECT 119.495 142.105 119.830 143.075 ;
        RECT 120.045 142.105 120.275 143.245 ;
        RECT 118.815 141.605 119.010 141.935 ;
        RECT 119.235 141.605 119.490 141.935 ;
        RECT 119.235 141.435 119.405 141.605 ;
        RECT 119.660 141.435 119.830 142.105 ;
        RECT 120.445 142.095 120.775 143.075 ;
        RECT 120.945 142.105 121.155 143.245 ;
        RECT 121.385 142.155 122.595 143.245 ;
        RECT 122.765 142.155 126.275 143.245 ;
        RECT 126.445 142.155 127.655 143.245 ;
        RECT 120.025 141.685 120.355 141.935 ;
        RECT 118.475 141.265 119.405 141.435 ;
        RECT 118.475 141.230 118.650 141.265 ;
        RECT 118.120 140.865 118.650 141.230 ;
        RECT 119.075 140.695 119.405 141.095 ;
        RECT 119.575 140.865 119.830 141.435 ;
        RECT 120.045 140.695 120.275 141.515 ;
        RECT 120.525 141.495 120.775 142.095 ;
        RECT 121.385 141.615 121.905 142.155 ;
        RECT 120.445 140.865 120.775 141.495 ;
        RECT 120.945 140.695 121.155 141.515 ;
        RECT 122.075 141.445 122.595 141.985 ;
        RECT 122.765 141.635 124.455 142.155 ;
        RECT 124.625 141.465 126.275 141.985 ;
        RECT 126.445 141.615 126.965 142.155 ;
        RECT 121.385 140.695 122.595 141.445 ;
        RECT 122.765 140.695 126.275 141.465 ;
        RECT 127.135 141.445 127.655 141.985 ;
        RECT 126.445 140.695 127.655 141.445 ;
        RECT 14.580 140.525 127.740 140.695 ;
        RECT 14.665 139.775 15.875 140.525 ;
        RECT 16.420 139.815 16.675 140.345 ;
        RECT 16.855 140.065 17.140 140.525 ;
        RECT 14.665 139.235 15.185 139.775 ;
        RECT 15.355 139.065 15.875 139.605 ;
        RECT 14.665 137.975 15.875 139.065 ;
        RECT 16.420 138.955 16.600 139.815 ;
        RECT 17.320 139.615 17.570 140.265 ;
        RECT 16.770 139.285 17.570 139.615 ;
        RECT 16.420 138.485 16.675 138.955 ;
        RECT 16.335 138.315 16.675 138.485 ;
        RECT 16.420 138.285 16.675 138.315 ;
        RECT 16.855 137.975 17.140 138.775 ;
        RECT 17.320 138.695 17.570 139.285 ;
        RECT 17.770 139.930 18.090 140.260 ;
        RECT 18.270 140.045 18.930 140.525 ;
        RECT 19.130 140.135 19.980 140.305 ;
        RECT 17.770 139.035 17.960 139.930 ;
        RECT 18.280 139.605 18.940 139.875 ;
        RECT 18.610 139.545 18.940 139.605 ;
        RECT 18.130 139.375 18.460 139.435 ;
        RECT 19.130 139.375 19.300 140.135 ;
        RECT 20.540 140.065 20.860 140.525 ;
        RECT 21.060 139.885 21.310 140.315 ;
        RECT 21.600 140.085 22.010 140.525 ;
        RECT 22.180 140.145 23.195 140.345 ;
        RECT 19.470 139.715 20.720 139.885 ;
        RECT 19.470 139.595 19.800 139.715 ;
        RECT 18.130 139.205 20.030 139.375 ;
        RECT 17.770 138.865 19.690 139.035 ;
        RECT 17.770 138.845 18.090 138.865 ;
        RECT 17.320 138.185 17.650 138.695 ;
        RECT 17.920 138.235 18.090 138.845 ;
        RECT 19.860 138.695 20.030 139.205 ;
        RECT 20.200 139.135 20.380 139.545 ;
        RECT 20.550 138.955 20.720 139.715 ;
        RECT 18.260 137.975 18.590 138.665 ;
        RECT 18.820 138.525 20.030 138.695 ;
        RECT 20.200 138.645 20.720 138.955 ;
        RECT 20.890 139.545 21.310 139.885 ;
        RECT 21.600 139.545 22.010 139.875 ;
        RECT 20.890 138.775 21.080 139.545 ;
        RECT 22.180 139.415 22.350 140.145 ;
        RECT 23.495 139.975 23.665 140.305 ;
        RECT 23.835 140.145 24.165 140.525 ;
        RECT 22.520 139.595 22.870 139.965 ;
        RECT 22.180 139.375 22.600 139.415 ;
        RECT 21.250 139.205 22.600 139.375 ;
        RECT 21.250 139.045 21.500 139.205 ;
        RECT 22.010 138.775 22.260 139.035 ;
        RECT 20.890 138.525 22.260 138.775 ;
        RECT 18.820 138.235 19.060 138.525 ;
        RECT 19.860 138.445 20.030 138.525 ;
        RECT 19.260 137.975 19.680 138.355 ;
        RECT 19.860 138.195 20.490 138.445 ;
        RECT 20.960 137.975 21.290 138.355 ;
        RECT 21.460 138.235 21.630 138.525 ;
        RECT 22.430 138.360 22.600 139.205 ;
        RECT 23.050 139.035 23.270 139.905 ;
        RECT 23.495 139.785 24.190 139.975 ;
        RECT 22.770 138.655 23.270 139.035 ;
        RECT 23.440 138.985 23.850 139.605 ;
        RECT 24.020 138.815 24.190 139.785 ;
        RECT 23.495 138.645 24.190 138.815 ;
        RECT 21.810 137.975 22.190 138.355 ;
        RECT 22.430 138.190 23.260 138.360 ;
        RECT 23.495 138.145 23.665 138.645 ;
        RECT 23.835 137.975 24.165 138.475 ;
        RECT 24.380 138.145 24.605 140.265 ;
        RECT 24.775 140.145 25.105 140.525 ;
        RECT 25.275 139.975 25.445 140.265 ;
        RECT 24.780 139.805 25.445 139.975 ;
        RECT 24.780 138.815 25.010 139.805 ;
        RECT 25.705 139.755 28.295 140.525 ;
        RECT 28.470 139.980 33.815 140.525 ;
        RECT 25.180 138.985 25.530 139.635 ;
        RECT 25.705 139.065 26.915 139.585 ;
        RECT 27.085 139.235 28.295 139.755 ;
        RECT 24.780 138.645 25.445 138.815 ;
        RECT 24.775 137.975 25.105 138.475 ;
        RECT 25.275 138.145 25.445 138.645 ;
        RECT 25.705 137.975 28.295 139.065 ;
        RECT 30.060 138.410 30.410 139.660 ;
        RECT 31.890 139.150 32.230 139.980 ;
        RECT 34.185 139.895 34.515 140.255 ;
        RECT 35.135 140.065 35.385 140.525 ;
        RECT 35.555 140.065 36.115 140.355 ;
        RECT 34.185 139.705 35.575 139.895 ;
        RECT 35.405 139.615 35.575 139.705 ;
        RECT 34.000 139.285 34.675 139.535 ;
        RECT 34.895 139.285 35.235 139.535 ;
        RECT 35.405 139.285 35.695 139.615 ;
        RECT 34.000 138.925 34.265 139.285 ;
        RECT 35.405 139.035 35.575 139.285 ;
        RECT 34.635 138.865 35.575 139.035 ;
        RECT 28.470 137.975 33.815 138.410 ;
        RECT 34.185 137.975 34.465 138.645 ;
        RECT 34.635 138.315 34.935 138.865 ;
        RECT 35.865 138.695 36.115 140.065 ;
        RECT 37.205 139.800 37.495 140.525 ;
        RECT 38.585 139.850 38.855 140.195 ;
        RECT 39.045 140.125 39.425 140.525 ;
        RECT 39.595 139.955 39.765 140.305 ;
        RECT 39.935 140.125 40.265 140.525 ;
        RECT 40.465 139.955 40.635 140.305 ;
        RECT 40.835 140.025 41.165 140.525 ;
        RECT 35.135 137.975 35.465 138.695 ;
        RECT 35.655 138.145 36.115 138.695 ;
        RECT 37.205 137.975 37.495 139.140 ;
        RECT 38.585 139.115 38.755 139.850 ;
        RECT 39.025 139.785 40.635 139.955 ;
        RECT 39.025 139.615 39.195 139.785 ;
        RECT 38.925 139.285 39.195 139.615 ;
        RECT 39.365 139.285 39.770 139.615 ;
        RECT 39.025 139.115 39.195 139.285 ;
        RECT 38.585 138.145 38.855 139.115 ;
        RECT 39.025 138.945 39.750 139.115 ;
        RECT 39.940 138.995 40.650 139.615 ;
        RECT 40.820 139.285 41.170 139.855 ;
        RECT 41.805 139.755 44.395 140.525 ;
        RECT 44.570 139.980 49.915 140.525 ;
        RECT 50.090 139.980 55.435 140.525 ;
        RECT 39.580 138.825 39.750 138.945 ;
        RECT 40.850 138.825 41.170 139.115 ;
        RECT 39.065 137.975 39.345 138.775 ;
        RECT 39.580 138.655 41.170 138.825 ;
        RECT 41.805 139.065 43.015 139.585 ;
        RECT 43.185 139.235 44.395 139.755 ;
        RECT 39.515 138.195 41.170 138.485 ;
        RECT 41.805 137.975 44.395 139.065 ;
        RECT 46.160 138.410 46.510 139.660 ;
        RECT 47.990 139.150 48.330 139.980 ;
        RECT 51.680 138.410 52.030 139.660 ;
        RECT 53.510 139.150 53.850 139.980 ;
        RECT 55.645 139.705 55.875 140.525 ;
        RECT 56.045 139.725 56.375 140.355 ;
        RECT 55.625 139.285 55.955 139.535 ;
        RECT 56.125 139.125 56.375 139.725 ;
        RECT 56.545 139.705 56.755 140.525 ;
        RECT 57.445 139.755 59.115 140.525 ;
        RECT 44.570 137.975 49.915 138.410 ;
        RECT 50.090 137.975 55.435 138.410 ;
        RECT 55.645 137.975 55.875 139.115 ;
        RECT 56.045 138.145 56.375 139.125 ;
        RECT 56.545 137.975 56.755 139.115 ;
        RECT 57.445 139.065 58.195 139.585 ;
        RECT 58.365 139.235 59.115 139.755 ;
        RECT 59.285 139.725 59.625 140.355 ;
        RECT 59.795 139.725 60.045 140.525 ;
        RECT 60.235 139.875 60.565 140.355 ;
        RECT 60.735 140.065 60.960 140.525 ;
        RECT 61.130 139.875 61.460 140.355 ;
        RECT 59.285 139.115 59.460 139.725 ;
        RECT 60.235 139.705 61.460 139.875 ;
        RECT 62.090 139.745 62.590 140.355 ;
        RECT 62.965 139.800 63.255 140.525 ;
        RECT 59.630 139.365 60.325 139.535 ;
        RECT 60.155 139.115 60.325 139.365 ;
        RECT 60.500 139.335 60.920 139.535 ;
        RECT 61.090 139.335 61.420 139.535 ;
        RECT 61.590 139.335 61.920 139.535 ;
        RECT 62.090 139.115 62.260 139.745 ;
        RECT 63.885 139.725 64.225 140.355 ;
        RECT 64.395 139.725 64.645 140.525 ;
        RECT 64.835 139.875 65.165 140.355 ;
        RECT 65.335 140.065 65.560 140.525 ;
        RECT 65.730 139.875 66.060 140.355 ;
        RECT 62.445 139.285 62.795 139.535 ;
        RECT 57.445 137.975 59.115 139.065 ;
        RECT 59.285 138.145 59.625 139.115 ;
        RECT 59.795 137.975 59.965 139.115 ;
        RECT 60.155 138.945 62.590 139.115 ;
        RECT 60.235 137.975 60.485 138.775 ;
        RECT 61.130 138.145 61.460 138.945 ;
        RECT 61.760 137.975 62.090 138.775 ;
        RECT 62.260 138.145 62.590 138.945 ;
        RECT 62.965 137.975 63.255 139.140 ;
        RECT 63.885 139.115 64.060 139.725 ;
        RECT 64.835 139.705 66.060 139.875 ;
        RECT 66.690 139.745 67.190 140.355 ;
        RECT 67.940 140.185 68.195 140.345 ;
        RECT 67.855 140.015 68.195 140.185 ;
        RECT 68.375 140.065 68.660 140.525 ;
        RECT 67.940 139.815 68.195 140.015 ;
        RECT 64.230 139.365 64.925 139.535 ;
        RECT 64.755 139.115 64.925 139.365 ;
        RECT 65.100 139.335 65.520 139.535 ;
        RECT 65.690 139.335 66.020 139.535 ;
        RECT 66.190 139.335 66.520 139.535 ;
        RECT 66.690 139.115 66.860 139.745 ;
        RECT 67.045 139.285 67.395 139.535 ;
        RECT 63.885 138.145 64.225 139.115 ;
        RECT 64.395 137.975 64.565 139.115 ;
        RECT 64.755 138.945 67.190 139.115 ;
        RECT 64.835 137.975 65.085 138.775 ;
        RECT 65.730 138.145 66.060 138.945 ;
        RECT 66.360 137.975 66.690 138.775 ;
        RECT 66.860 138.145 67.190 138.945 ;
        RECT 67.940 138.955 68.120 139.815 ;
        RECT 68.840 139.615 69.090 140.265 ;
        RECT 68.290 139.285 69.090 139.615 ;
        RECT 67.940 138.285 68.195 138.955 ;
        RECT 68.375 137.975 68.660 138.775 ;
        RECT 68.840 138.695 69.090 139.285 ;
        RECT 69.290 139.930 69.610 140.260 ;
        RECT 69.790 140.045 70.450 140.525 ;
        RECT 70.650 140.135 71.500 140.305 ;
        RECT 69.290 139.035 69.480 139.930 ;
        RECT 69.800 139.605 70.460 139.875 ;
        RECT 70.130 139.545 70.460 139.605 ;
        RECT 69.650 139.375 69.980 139.435 ;
        RECT 70.650 139.375 70.820 140.135 ;
        RECT 72.060 140.065 72.380 140.525 ;
        RECT 72.580 139.885 72.830 140.315 ;
        RECT 73.120 140.085 73.530 140.525 ;
        RECT 73.700 140.145 74.715 140.345 ;
        RECT 70.990 139.715 72.240 139.885 ;
        RECT 70.990 139.595 71.320 139.715 ;
        RECT 69.650 139.205 71.550 139.375 ;
        RECT 69.290 138.865 71.210 139.035 ;
        RECT 69.290 138.845 69.610 138.865 ;
        RECT 68.840 138.185 69.170 138.695 ;
        RECT 69.440 138.235 69.610 138.845 ;
        RECT 71.380 138.695 71.550 139.205 ;
        RECT 71.720 139.135 71.900 139.545 ;
        RECT 72.070 138.955 72.240 139.715 ;
        RECT 69.780 137.975 70.110 138.665 ;
        RECT 70.340 138.525 71.550 138.695 ;
        RECT 71.720 138.645 72.240 138.955 ;
        RECT 72.410 139.545 72.830 139.885 ;
        RECT 73.120 139.545 73.530 139.875 ;
        RECT 72.410 138.775 72.600 139.545 ;
        RECT 73.700 139.415 73.870 140.145 ;
        RECT 75.015 139.975 75.185 140.305 ;
        RECT 75.355 140.145 75.685 140.525 ;
        RECT 74.040 139.595 74.390 139.965 ;
        RECT 73.700 139.375 74.120 139.415 ;
        RECT 72.770 139.205 74.120 139.375 ;
        RECT 72.770 139.045 73.020 139.205 ;
        RECT 73.530 138.775 73.780 139.035 ;
        RECT 72.410 138.525 73.780 138.775 ;
        RECT 70.340 138.235 70.580 138.525 ;
        RECT 71.380 138.445 71.550 138.525 ;
        RECT 70.780 137.975 71.200 138.355 ;
        RECT 71.380 138.195 72.010 138.445 ;
        RECT 72.480 137.975 72.810 138.355 ;
        RECT 72.980 138.235 73.150 138.525 ;
        RECT 73.950 138.360 74.120 139.205 ;
        RECT 74.570 139.035 74.790 139.905 ;
        RECT 75.015 139.785 75.710 139.975 ;
        RECT 74.290 138.655 74.790 139.035 ;
        RECT 74.960 138.985 75.370 139.605 ;
        RECT 75.540 138.815 75.710 139.785 ;
        RECT 75.015 138.645 75.710 138.815 ;
        RECT 73.330 137.975 73.710 138.355 ;
        RECT 73.950 138.190 74.780 138.360 ;
        RECT 75.015 138.145 75.185 138.645 ;
        RECT 75.355 137.975 75.685 138.475 ;
        RECT 75.900 138.145 76.125 140.265 ;
        RECT 76.295 140.145 76.625 140.525 ;
        RECT 76.795 139.975 76.965 140.265 ;
        RECT 76.300 139.805 76.965 139.975 ;
        RECT 76.300 138.815 76.530 139.805 ;
        RECT 77.685 139.755 79.355 140.525 ;
        RECT 76.700 138.985 77.050 139.635 ;
        RECT 77.685 139.065 78.435 139.585 ;
        RECT 78.605 139.235 79.355 139.755 ;
        RECT 79.525 139.725 79.865 140.355 ;
        RECT 80.035 139.725 80.285 140.525 ;
        RECT 80.475 139.875 80.805 140.355 ;
        RECT 80.975 140.065 81.200 140.525 ;
        RECT 81.370 139.875 81.700 140.355 ;
        RECT 79.525 139.115 79.700 139.725 ;
        RECT 80.475 139.705 81.700 139.875 ;
        RECT 82.330 139.745 82.830 140.355 ;
        RECT 83.205 139.775 84.415 140.525 ;
        RECT 79.870 139.365 80.565 139.535 ;
        RECT 80.395 139.115 80.565 139.365 ;
        RECT 80.740 139.335 81.160 139.535 ;
        RECT 81.330 139.335 81.660 139.535 ;
        RECT 81.830 139.335 82.160 139.535 ;
        RECT 82.330 139.115 82.500 139.745 ;
        RECT 82.685 139.285 83.035 139.535 ;
        RECT 76.300 138.645 76.965 138.815 ;
        RECT 76.295 137.975 76.625 138.475 ;
        RECT 76.795 138.145 76.965 138.645 ;
        RECT 77.685 137.975 79.355 139.065 ;
        RECT 79.525 138.145 79.865 139.115 ;
        RECT 80.035 137.975 80.205 139.115 ;
        RECT 80.395 138.945 82.830 139.115 ;
        RECT 80.475 137.975 80.725 138.775 ;
        RECT 81.370 138.145 81.700 138.945 ;
        RECT 82.000 137.975 82.330 138.775 ;
        RECT 82.500 138.145 82.830 138.945 ;
        RECT 83.205 139.065 83.725 139.605 ;
        RECT 83.895 139.235 84.415 139.775 ;
        RECT 84.860 139.715 85.105 140.320 ;
        RECT 85.325 139.990 85.835 140.525 ;
        RECT 84.585 139.545 85.815 139.715 ;
        RECT 83.205 137.975 84.415 139.065 ;
        RECT 84.585 138.735 84.925 139.545 ;
        RECT 85.095 138.980 85.845 139.170 ;
        RECT 84.585 138.325 85.100 138.735 ;
        RECT 85.335 137.975 85.505 138.735 ;
        RECT 85.675 138.315 85.845 138.980 ;
        RECT 86.015 138.995 86.205 140.355 ;
        RECT 86.375 139.505 86.650 140.355 ;
        RECT 86.840 139.990 87.370 140.355 ;
        RECT 87.795 140.125 88.125 140.525 ;
        RECT 87.195 139.955 87.370 139.990 ;
        RECT 86.375 139.335 86.655 139.505 ;
        RECT 86.375 139.195 86.650 139.335 ;
        RECT 86.855 138.995 87.025 139.795 ;
        RECT 86.015 138.825 87.025 138.995 ;
        RECT 87.195 139.785 88.125 139.955 ;
        RECT 88.295 139.785 88.550 140.355 ;
        RECT 88.725 139.800 89.015 140.525 ;
        RECT 89.275 139.975 89.445 140.355 ;
        RECT 89.625 140.145 89.955 140.525 ;
        RECT 89.275 139.805 89.940 139.975 ;
        RECT 90.135 139.850 90.395 140.355 ;
        RECT 87.195 138.655 87.365 139.785 ;
        RECT 87.955 139.615 88.125 139.785 ;
        RECT 86.240 138.485 87.365 138.655 ;
        RECT 87.535 139.285 87.730 139.615 ;
        RECT 87.955 139.285 88.210 139.615 ;
        RECT 87.535 138.315 87.705 139.285 ;
        RECT 88.380 139.115 88.550 139.785 ;
        RECT 89.205 139.255 89.535 139.625 ;
        RECT 89.770 139.550 89.940 139.805 ;
        RECT 89.770 139.220 90.055 139.550 ;
        RECT 85.675 138.145 87.705 138.315 ;
        RECT 87.875 137.975 88.045 139.115 ;
        RECT 88.215 138.145 88.550 139.115 ;
        RECT 88.725 137.975 89.015 139.140 ;
        RECT 89.770 139.075 89.940 139.220 ;
        RECT 89.275 138.905 89.940 139.075 ;
        RECT 90.225 139.050 90.395 139.850 ;
        RECT 90.565 139.755 92.235 140.525 ;
        RECT 92.410 139.980 97.755 140.525 ;
        RECT 89.275 138.145 89.445 138.905 ;
        RECT 89.625 137.975 89.955 138.735 ;
        RECT 90.125 138.145 90.395 139.050 ;
        RECT 90.565 139.065 91.315 139.585 ;
        RECT 91.485 139.235 92.235 139.755 ;
        RECT 90.565 137.975 92.235 139.065 ;
        RECT 94.000 138.410 94.350 139.660 ;
        RECT 95.830 139.150 96.170 139.980 ;
        RECT 98.300 139.815 98.555 140.345 ;
        RECT 98.735 140.065 99.020 140.525 ;
        RECT 98.300 139.165 98.480 139.815 ;
        RECT 99.200 139.615 99.450 140.265 ;
        RECT 98.650 139.285 99.450 139.615 ;
        RECT 98.215 138.995 98.480 139.165 ;
        RECT 98.300 138.955 98.480 138.995 ;
        RECT 92.410 137.975 97.755 138.410 ;
        RECT 98.300 138.285 98.555 138.955 ;
        RECT 98.735 137.975 99.020 138.775 ;
        RECT 99.200 138.695 99.450 139.285 ;
        RECT 99.650 139.930 99.970 140.260 ;
        RECT 100.150 140.045 100.810 140.525 ;
        RECT 101.010 140.135 101.860 140.305 ;
        RECT 99.650 139.035 99.840 139.930 ;
        RECT 100.160 139.605 100.820 139.875 ;
        RECT 100.490 139.545 100.820 139.605 ;
        RECT 100.010 139.375 100.340 139.435 ;
        RECT 101.010 139.375 101.180 140.135 ;
        RECT 102.420 140.065 102.740 140.525 ;
        RECT 102.940 139.885 103.190 140.315 ;
        RECT 103.480 140.085 103.890 140.525 ;
        RECT 104.060 140.145 105.075 140.345 ;
        RECT 101.350 139.715 102.600 139.885 ;
        RECT 101.350 139.595 101.680 139.715 ;
        RECT 100.010 139.205 101.910 139.375 ;
        RECT 99.650 138.865 101.570 139.035 ;
        RECT 99.650 138.845 99.970 138.865 ;
        RECT 99.200 138.185 99.530 138.695 ;
        RECT 99.800 138.235 99.970 138.845 ;
        RECT 101.740 138.695 101.910 139.205 ;
        RECT 102.080 139.135 102.260 139.545 ;
        RECT 102.430 138.955 102.600 139.715 ;
        RECT 100.140 137.975 100.470 138.665 ;
        RECT 100.700 138.525 101.910 138.695 ;
        RECT 102.080 138.645 102.600 138.955 ;
        RECT 102.770 139.545 103.190 139.885 ;
        RECT 103.480 139.545 103.890 139.875 ;
        RECT 102.770 138.775 102.960 139.545 ;
        RECT 104.060 139.415 104.230 140.145 ;
        RECT 105.375 139.975 105.545 140.305 ;
        RECT 105.715 140.145 106.045 140.525 ;
        RECT 104.400 139.595 104.750 139.965 ;
        RECT 104.060 139.375 104.480 139.415 ;
        RECT 103.130 139.205 104.480 139.375 ;
        RECT 103.130 139.045 103.380 139.205 ;
        RECT 103.890 138.775 104.140 139.035 ;
        RECT 102.770 138.525 104.140 138.775 ;
        RECT 100.700 138.235 100.940 138.525 ;
        RECT 101.740 138.445 101.910 138.525 ;
        RECT 101.140 137.975 101.560 138.355 ;
        RECT 101.740 138.195 102.370 138.445 ;
        RECT 102.840 137.975 103.170 138.355 ;
        RECT 103.340 138.235 103.510 138.525 ;
        RECT 104.310 138.360 104.480 139.205 ;
        RECT 104.930 139.035 105.150 139.905 ;
        RECT 105.375 139.785 106.070 139.975 ;
        RECT 104.650 138.655 105.150 139.035 ;
        RECT 105.320 138.985 105.730 139.605 ;
        RECT 105.900 138.815 106.070 139.785 ;
        RECT 105.375 138.645 106.070 138.815 ;
        RECT 103.690 137.975 104.070 138.355 ;
        RECT 104.310 138.190 105.140 138.360 ;
        RECT 105.375 138.145 105.545 138.645 ;
        RECT 105.715 137.975 106.045 138.475 ;
        RECT 106.260 138.145 106.485 140.265 ;
        RECT 106.655 140.145 106.985 140.525 ;
        RECT 107.155 139.975 107.325 140.265 ;
        RECT 106.660 139.805 107.325 139.975 ;
        RECT 106.660 138.815 106.890 139.805 ;
        RECT 108.045 139.755 109.715 140.525 ;
        RECT 107.060 138.985 107.410 139.635 ;
        RECT 108.045 139.065 108.795 139.585 ;
        RECT 108.965 139.235 109.715 139.755 ;
        RECT 110.090 139.745 110.590 140.355 ;
        RECT 109.885 139.285 110.235 139.535 ;
        RECT 110.420 139.115 110.590 139.745 ;
        RECT 111.220 139.875 111.550 140.355 ;
        RECT 111.720 140.065 111.945 140.525 ;
        RECT 112.115 139.875 112.445 140.355 ;
        RECT 111.220 139.705 112.445 139.875 ;
        RECT 112.635 139.725 112.885 140.525 ;
        RECT 113.055 139.725 113.395 140.355 ;
        RECT 114.485 139.800 114.775 140.525 ;
        RECT 113.165 139.675 113.395 139.725 ;
        RECT 115.445 139.705 115.675 140.525 ;
        RECT 115.845 139.725 116.175 140.355 ;
        RECT 110.760 139.335 111.090 139.535 ;
        RECT 111.260 139.335 111.590 139.535 ;
        RECT 111.760 139.335 112.180 139.535 ;
        RECT 112.355 139.365 113.050 139.535 ;
        RECT 112.355 139.115 112.525 139.365 ;
        RECT 113.220 139.115 113.395 139.675 ;
        RECT 115.425 139.285 115.755 139.535 ;
        RECT 106.660 138.645 107.325 138.815 ;
        RECT 106.655 137.975 106.985 138.475 ;
        RECT 107.155 138.145 107.325 138.645 ;
        RECT 108.045 137.975 109.715 139.065 ;
        RECT 110.090 138.945 112.525 139.115 ;
        RECT 110.090 138.145 110.420 138.945 ;
        RECT 110.590 137.975 110.920 138.775 ;
        RECT 111.220 138.145 111.550 138.945 ;
        RECT 112.195 137.975 112.445 138.775 ;
        RECT 112.715 137.975 112.885 139.115 ;
        RECT 113.055 138.145 113.395 139.115 ;
        RECT 114.485 137.975 114.775 139.140 ;
        RECT 115.925 139.125 116.175 139.725 ;
        RECT 116.345 139.705 116.555 140.525 ;
        RECT 117.160 139.845 117.415 140.345 ;
        RECT 117.595 140.065 117.880 140.525 ;
        RECT 117.075 139.815 117.415 139.845 ;
        RECT 117.075 139.675 117.340 139.815 ;
        RECT 115.445 137.975 115.675 139.115 ;
        RECT 115.845 138.145 116.175 139.125 ;
        RECT 116.345 137.975 116.555 139.115 ;
        RECT 117.160 138.955 117.340 139.675 ;
        RECT 118.060 139.615 118.310 140.265 ;
        RECT 117.510 139.285 118.310 139.615 ;
        RECT 117.160 138.285 117.415 138.955 ;
        RECT 117.595 137.975 117.880 138.775 ;
        RECT 118.060 138.695 118.310 139.285 ;
        RECT 118.510 139.930 118.830 140.260 ;
        RECT 119.010 140.045 119.670 140.525 ;
        RECT 119.870 140.135 120.720 140.305 ;
        RECT 118.510 139.035 118.700 139.930 ;
        RECT 119.020 139.605 119.680 139.875 ;
        RECT 119.350 139.545 119.680 139.605 ;
        RECT 118.870 139.375 119.200 139.435 ;
        RECT 119.870 139.375 120.040 140.135 ;
        RECT 121.280 140.065 121.600 140.525 ;
        RECT 121.800 139.885 122.050 140.315 ;
        RECT 122.340 140.085 122.750 140.525 ;
        RECT 122.920 140.145 123.935 140.345 ;
        RECT 120.210 139.715 121.460 139.885 ;
        RECT 120.210 139.595 120.540 139.715 ;
        RECT 118.870 139.205 120.770 139.375 ;
        RECT 118.510 138.865 120.430 139.035 ;
        RECT 118.510 138.845 118.830 138.865 ;
        RECT 118.060 138.185 118.390 138.695 ;
        RECT 118.660 138.235 118.830 138.845 ;
        RECT 120.600 138.695 120.770 139.205 ;
        RECT 120.940 139.135 121.120 139.545 ;
        RECT 121.290 138.955 121.460 139.715 ;
        RECT 119.000 137.975 119.330 138.665 ;
        RECT 119.560 138.525 120.770 138.695 ;
        RECT 120.940 138.645 121.460 138.955 ;
        RECT 121.630 139.545 122.050 139.885 ;
        RECT 122.340 139.545 122.750 139.875 ;
        RECT 121.630 138.775 121.820 139.545 ;
        RECT 122.920 139.415 123.090 140.145 ;
        RECT 124.235 139.975 124.405 140.305 ;
        RECT 124.575 140.145 124.905 140.525 ;
        RECT 123.260 139.595 123.610 139.965 ;
        RECT 122.920 139.375 123.340 139.415 ;
        RECT 121.990 139.205 123.340 139.375 ;
        RECT 121.990 139.045 122.240 139.205 ;
        RECT 122.750 138.775 123.000 139.035 ;
        RECT 121.630 138.525 123.000 138.775 ;
        RECT 119.560 138.235 119.800 138.525 ;
        RECT 120.600 138.445 120.770 138.525 ;
        RECT 120.000 137.975 120.420 138.355 ;
        RECT 120.600 138.195 121.230 138.445 ;
        RECT 121.700 137.975 122.030 138.355 ;
        RECT 122.200 138.235 122.370 138.525 ;
        RECT 123.170 138.360 123.340 139.205 ;
        RECT 123.790 139.035 124.010 139.905 ;
        RECT 124.235 139.785 124.930 139.975 ;
        RECT 123.510 138.655 124.010 139.035 ;
        RECT 124.180 138.985 124.590 139.605 ;
        RECT 124.760 138.815 124.930 139.785 ;
        RECT 124.235 138.645 124.930 138.815 ;
        RECT 122.550 137.975 122.930 138.355 ;
        RECT 123.170 138.190 124.000 138.360 ;
        RECT 124.235 138.145 124.405 138.645 ;
        RECT 124.575 137.975 124.905 138.475 ;
        RECT 125.120 138.145 125.345 140.265 ;
        RECT 125.515 140.145 125.845 140.525 ;
        RECT 126.015 139.975 126.185 140.265 ;
        RECT 125.520 139.805 126.185 139.975 ;
        RECT 125.520 138.815 125.750 139.805 ;
        RECT 126.445 139.775 127.655 140.525 ;
        RECT 125.920 138.985 126.270 139.635 ;
        RECT 126.445 139.065 126.965 139.605 ;
        RECT 127.135 139.235 127.655 139.775 ;
        RECT 125.520 138.645 126.185 138.815 ;
        RECT 125.515 137.975 125.845 138.475 ;
        RECT 126.015 138.145 126.185 138.645 ;
        RECT 126.445 137.975 127.655 139.065 ;
        RECT 14.580 137.805 127.740 137.975 ;
        RECT 14.665 136.715 15.875 137.805 ;
        RECT 14.665 136.005 15.185 136.545 ;
        RECT 15.355 136.175 15.875 136.715 ;
        RECT 16.505 136.715 20.015 137.805 ;
        RECT 16.505 136.195 18.195 136.715 ;
        RECT 20.190 136.665 20.525 137.635 ;
        RECT 20.695 136.665 20.865 137.805 ;
        RECT 21.035 137.465 23.065 137.635 ;
        RECT 18.365 136.025 20.015 136.545 ;
        RECT 14.665 135.255 15.875 136.005 ;
        RECT 16.505 135.255 20.015 136.025 ;
        RECT 20.190 135.995 20.360 136.665 ;
        RECT 21.035 136.495 21.205 137.465 ;
        RECT 20.530 136.165 20.785 136.495 ;
        RECT 21.010 136.165 21.205 136.495 ;
        RECT 21.375 137.125 22.500 137.295 ;
        RECT 20.615 135.995 20.785 136.165 ;
        RECT 21.375 135.995 21.545 137.125 ;
        RECT 20.190 135.425 20.445 135.995 ;
        RECT 20.615 135.825 21.545 135.995 ;
        RECT 21.715 136.785 22.725 136.955 ;
        RECT 21.715 135.985 21.885 136.785 ;
        RECT 22.090 136.445 22.365 136.585 ;
        RECT 22.085 136.275 22.365 136.445 ;
        RECT 21.370 135.790 21.545 135.825 ;
        RECT 20.615 135.255 20.945 135.655 ;
        RECT 21.370 135.425 21.900 135.790 ;
        RECT 22.090 135.425 22.365 136.275 ;
        RECT 22.535 135.425 22.725 136.785 ;
        RECT 22.895 136.800 23.065 137.465 ;
        RECT 23.235 137.045 23.405 137.805 ;
        RECT 23.640 137.045 24.155 137.455 ;
        RECT 22.895 136.610 23.645 136.800 ;
        RECT 23.815 136.235 24.155 137.045 ;
        RECT 24.325 136.640 24.615 137.805 ;
        RECT 24.785 136.715 28.295 137.805 ;
        RECT 22.925 136.065 24.155 136.235 ;
        RECT 24.785 136.195 26.475 136.715 ;
        RECT 28.470 136.665 28.805 137.635 ;
        RECT 28.975 136.665 29.145 137.805 ;
        RECT 29.315 137.465 31.345 137.635 ;
        RECT 22.905 135.255 23.415 135.790 ;
        RECT 23.635 135.460 23.880 136.065 ;
        RECT 26.645 136.025 28.295 136.545 ;
        RECT 24.325 135.255 24.615 135.980 ;
        RECT 24.785 135.255 28.295 136.025 ;
        RECT 28.470 135.995 28.640 136.665 ;
        RECT 29.315 136.495 29.485 137.465 ;
        RECT 28.810 136.165 29.065 136.495 ;
        RECT 29.290 136.165 29.485 136.495 ;
        RECT 29.655 137.125 30.780 137.295 ;
        RECT 28.895 135.995 29.065 136.165 ;
        RECT 29.655 135.995 29.825 137.125 ;
        RECT 28.470 135.425 28.725 135.995 ;
        RECT 28.895 135.825 29.825 135.995 ;
        RECT 29.995 136.785 31.005 136.955 ;
        RECT 29.995 135.985 30.165 136.785 ;
        RECT 30.370 136.105 30.645 136.585 ;
        RECT 30.365 135.935 30.645 136.105 ;
        RECT 29.650 135.790 29.825 135.825 ;
        RECT 28.895 135.255 29.225 135.655 ;
        RECT 29.650 135.425 30.180 135.790 ;
        RECT 30.370 135.425 30.645 135.935 ;
        RECT 30.815 135.425 31.005 136.785 ;
        RECT 31.175 136.800 31.345 137.465 ;
        RECT 31.515 137.045 31.685 137.805 ;
        RECT 31.920 137.045 32.435 137.455 ;
        RECT 32.805 137.135 33.085 137.805 ;
        RECT 31.175 136.610 31.925 136.800 ;
        RECT 32.095 136.235 32.435 137.045 ;
        RECT 33.255 136.915 33.555 137.465 ;
        RECT 33.755 137.085 34.085 137.805 ;
        RECT 34.275 137.085 34.735 137.635 ;
        RECT 32.620 136.495 32.885 136.855 ;
        RECT 33.255 136.745 34.195 136.915 ;
        RECT 34.025 136.495 34.195 136.745 ;
        RECT 32.620 136.245 33.295 136.495 ;
        RECT 33.515 136.245 33.855 136.495 ;
        RECT 31.205 136.065 32.435 136.235 ;
        RECT 34.025 136.165 34.315 136.495 ;
        RECT 34.025 136.075 34.195 136.165 ;
        RECT 31.185 135.255 31.695 135.790 ;
        RECT 31.915 135.460 32.160 136.065 ;
        RECT 32.805 135.885 34.195 136.075 ;
        RECT 32.805 135.525 33.135 135.885 ;
        RECT 34.485 135.715 34.735 137.085 ;
        RECT 33.755 135.255 34.005 135.715 ;
        RECT 34.175 135.425 34.735 135.715 ;
        RECT 34.905 136.665 35.175 137.635 ;
        RECT 35.385 137.005 35.665 137.805 ;
        RECT 35.835 137.295 37.490 137.585 ;
        RECT 35.900 136.955 37.490 137.125 ;
        RECT 35.900 136.835 36.070 136.955 ;
        RECT 35.345 136.665 36.070 136.835 ;
        RECT 34.905 135.930 35.075 136.665 ;
        RECT 35.345 136.495 35.515 136.665 ;
        RECT 35.245 136.165 35.515 136.495 ;
        RECT 35.685 136.165 36.090 136.495 ;
        RECT 36.260 136.165 36.970 136.785 ;
        RECT 37.170 136.665 37.490 136.955 ;
        RECT 37.665 136.665 37.935 137.635 ;
        RECT 38.145 137.005 38.425 137.805 ;
        RECT 38.595 137.295 40.250 137.585 ;
        RECT 38.660 136.955 40.250 137.125 ;
        RECT 38.660 136.835 38.830 136.955 ;
        RECT 38.105 136.665 38.830 136.835 ;
        RECT 35.345 135.995 35.515 136.165 ;
        RECT 34.905 135.585 35.175 135.930 ;
        RECT 35.345 135.825 36.955 135.995 ;
        RECT 37.140 135.925 37.490 136.495 ;
        RECT 37.665 135.930 37.835 136.665 ;
        RECT 38.105 136.495 38.275 136.665 ;
        RECT 38.005 136.165 38.275 136.495 ;
        RECT 38.445 136.165 38.850 136.495 ;
        RECT 39.020 136.165 39.730 136.785 ;
        RECT 39.930 136.665 40.250 136.955 ;
        RECT 40.885 136.715 43.475 137.805 ;
        RECT 38.105 135.995 38.275 136.165 ;
        RECT 35.365 135.255 35.745 135.655 ;
        RECT 35.915 135.475 36.085 135.825 ;
        RECT 36.255 135.255 36.585 135.655 ;
        RECT 36.785 135.475 36.955 135.825 ;
        RECT 37.155 135.255 37.485 135.755 ;
        RECT 37.665 135.585 37.935 135.930 ;
        RECT 38.105 135.825 39.715 135.995 ;
        RECT 39.900 135.925 40.250 136.495 ;
        RECT 40.885 136.195 42.095 136.715 ;
        RECT 43.645 136.665 43.915 137.635 ;
        RECT 44.125 137.005 44.405 137.805 ;
        RECT 44.575 137.295 46.230 137.585 ;
        RECT 44.640 136.955 46.230 137.125 ;
        RECT 44.640 136.835 44.810 136.955 ;
        RECT 44.085 136.665 44.810 136.835 ;
        RECT 42.265 136.025 43.475 136.545 ;
        RECT 38.125 135.255 38.505 135.655 ;
        RECT 38.675 135.475 38.845 135.825 ;
        RECT 39.015 135.255 39.345 135.655 ;
        RECT 39.545 135.475 39.715 135.825 ;
        RECT 39.915 135.255 40.245 135.755 ;
        RECT 40.885 135.255 43.475 136.025 ;
        RECT 43.645 135.930 43.815 136.665 ;
        RECT 44.085 136.495 44.255 136.665 ;
        RECT 45.000 136.615 45.715 136.785 ;
        RECT 45.910 136.665 46.230 136.955 ;
        RECT 46.405 136.665 46.745 137.635 ;
        RECT 46.915 136.665 47.085 137.805 ;
        RECT 47.355 137.005 47.605 137.805 ;
        RECT 48.250 136.835 48.580 137.635 ;
        RECT 48.880 137.005 49.210 137.805 ;
        RECT 49.380 136.835 49.710 137.635 ;
        RECT 47.275 136.665 49.710 136.835 ;
        RECT 43.985 136.165 44.255 136.495 ;
        RECT 44.425 136.165 44.830 136.495 ;
        RECT 45.000 136.165 45.710 136.615 ;
        RECT 44.085 135.995 44.255 136.165 ;
        RECT 43.645 135.585 43.915 135.930 ;
        RECT 44.085 135.825 45.695 135.995 ;
        RECT 45.880 135.925 46.230 136.495 ;
        RECT 46.405 136.105 46.580 136.665 ;
        RECT 47.275 136.415 47.445 136.665 ;
        RECT 46.750 136.245 47.445 136.415 ;
        RECT 47.620 136.245 48.040 136.445 ;
        RECT 48.210 136.245 48.540 136.445 ;
        RECT 48.710 136.245 49.040 136.445 ;
        RECT 46.405 136.055 46.635 136.105 ;
        RECT 44.105 135.255 44.485 135.655 ;
        RECT 44.655 135.475 44.825 135.825 ;
        RECT 44.995 135.255 45.325 135.655 ;
        RECT 45.525 135.475 45.695 135.825 ;
        RECT 45.895 135.255 46.225 135.755 ;
        RECT 46.405 135.425 46.745 136.055 ;
        RECT 46.915 135.255 47.165 136.055 ;
        RECT 47.355 135.905 48.580 136.075 ;
        RECT 47.355 135.425 47.685 135.905 ;
        RECT 47.855 135.255 48.080 135.715 ;
        RECT 48.250 135.425 48.580 135.905 ;
        RECT 49.210 136.035 49.380 136.665 ;
        RECT 50.085 136.640 50.375 137.805 ;
        RECT 50.545 136.715 53.135 137.805 ;
        RECT 53.305 137.045 53.820 137.455 ;
        RECT 54.055 137.045 54.225 137.805 ;
        RECT 54.395 137.465 56.425 137.635 ;
        RECT 49.565 136.245 49.915 136.495 ;
        RECT 50.545 136.195 51.755 136.715 ;
        RECT 49.210 135.425 49.710 136.035 ;
        RECT 51.925 136.025 53.135 136.545 ;
        RECT 53.305 136.235 53.645 137.045 ;
        RECT 54.395 136.800 54.565 137.465 ;
        RECT 54.960 137.125 56.085 137.295 ;
        RECT 53.815 136.610 54.565 136.800 ;
        RECT 54.735 136.785 55.745 136.955 ;
        RECT 53.305 136.065 54.535 136.235 ;
        RECT 50.085 135.255 50.375 135.980 ;
        RECT 50.545 135.255 53.135 136.025 ;
        RECT 53.580 135.460 53.825 136.065 ;
        RECT 54.045 135.255 54.555 135.790 ;
        RECT 54.735 135.425 54.925 136.785 ;
        RECT 55.095 136.445 55.370 136.585 ;
        RECT 55.095 136.275 55.375 136.445 ;
        RECT 55.095 135.425 55.370 136.275 ;
        RECT 55.575 135.985 55.745 136.785 ;
        RECT 55.915 135.995 56.085 137.125 ;
        RECT 56.255 136.495 56.425 137.465 ;
        RECT 56.595 136.665 56.765 137.805 ;
        RECT 56.935 136.665 57.270 137.635 ;
        RECT 57.995 136.875 58.165 137.635 ;
        RECT 58.345 137.045 58.675 137.805 ;
        RECT 57.995 136.705 58.660 136.875 ;
        RECT 58.845 136.730 59.115 137.635 ;
        RECT 56.255 136.165 56.450 136.495 ;
        RECT 56.675 136.165 56.930 136.495 ;
        RECT 56.675 135.995 56.845 136.165 ;
        RECT 57.100 135.995 57.270 136.665 ;
        RECT 58.490 136.560 58.660 136.705 ;
        RECT 57.925 136.155 58.255 136.525 ;
        RECT 58.490 136.230 58.775 136.560 ;
        RECT 55.915 135.825 56.845 135.995 ;
        RECT 55.915 135.790 56.090 135.825 ;
        RECT 55.560 135.425 56.090 135.790 ;
        RECT 56.515 135.255 56.845 135.655 ;
        RECT 57.015 135.425 57.270 135.995 ;
        RECT 58.490 135.975 58.660 136.230 ;
        RECT 57.995 135.805 58.660 135.975 ;
        RECT 58.945 135.930 59.115 136.730 ;
        RECT 59.285 136.715 60.955 137.805 ;
        RECT 59.285 136.195 60.035 136.715 ;
        RECT 61.125 136.665 61.465 137.635 ;
        RECT 61.635 136.665 61.805 137.805 ;
        RECT 62.075 137.005 62.325 137.805 ;
        RECT 62.970 136.835 63.300 137.635 ;
        RECT 63.600 137.005 63.930 137.805 ;
        RECT 64.100 136.835 64.430 137.635 ;
        RECT 64.920 137.175 65.205 137.635 ;
        RECT 65.375 137.345 65.645 137.805 ;
        RECT 64.920 136.955 65.875 137.175 ;
        RECT 61.995 136.665 64.430 136.835 ;
        RECT 60.205 136.025 60.955 136.545 ;
        RECT 57.995 135.425 58.165 135.805 ;
        RECT 58.345 135.255 58.675 135.635 ;
        RECT 58.855 135.425 59.115 135.930 ;
        RECT 59.285 135.255 60.955 136.025 ;
        RECT 61.125 136.055 61.300 136.665 ;
        RECT 61.995 136.415 62.165 136.665 ;
        RECT 61.470 136.245 62.165 136.415 ;
        RECT 62.340 136.245 62.760 136.445 ;
        RECT 62.930 136.245 63.260 136.445 ;
        RECT 63.430 136.245 63.760 136.445 ;
        RECT 61.125 135.425 61.465 136.055 ;
        RECT 61.635 135.255 61.885 136.055 ;
        RECT 62.075 135.905 63.300 136.075 ;
        RECT 62.075 135.425 62.405 135.905 ;
        RECT 62.575 135.255 62.800 135.715 ;
        RECT 62.970 135.425 63.300 135.905 ;
        RECT 63.930 136.035 64.100 136.665 ;
        RECT 64.285 136.245 64.635 136.495 ;
        RECT 64.805 136.225 65.495 136.785 ;
        RECT 65.665 136.055 65.875 136.955 ;
        RECT 63.930 135.425 64.430 136.035 ;
        RECT 64.920 135.885 65.875 136.055 ;
        RECT 66.045 136.785 66.445 137.635 ;
        RECT 66.635 137.175 66.915 137.635 ;
        RECT 67.435 137.345 67.760 137.805 ;
        RECT 66.635 136.955 67.760 137.175 ;
        RECT 66.045 136.225 67.140 136.785 ;
        RECT 67.310 136.495 67.760 136.955 ;
        RECT 67.930 136.665 68.315 137.635 ;
        RECT 64.920 135.425 65.205 135.885 ;
        RECT 65.375 135.255 65.645 135.715 ;
        RECT 66.045 135.425 66.445 136.225 ;
        RECT 67.310 136.165 67.865 136.495 ;
        RECT 67.310 136.055 67.760 136.165 ;
        RECT 66.635 135.885 67.760 136.055 ;
        RECT 68.035 135.995 68.315 136.665 ;
        RECT 68.490 137.415 68.825 137.635 ;
        RECT 69.830 137.425 70.185 137.805 ;
        RECT 68.490 136.795 68.745 137.415 ;
        RECT 68.995 137.255 69.225 137.295 ;
        RECT 70.355 137.255 70.605 137.635 ;
        RECT 68.995 137.055 70.605 137.255 ;
        RECT 68.995 136.965 69.180 137.055 ;
        RECT 69.770 137.045 70.605 137.055 ;
        RECT 70.855 137.025 71.105 137.805 ;
        RECT 71.275 136.955 71.535 137.635 ;
        RECT 69.335 136.855 69.665 136.885 ;
        RECT 69.335 136.795 71.135 136.855 ;
        RECT 68.490 136.685 71.195 136.795 ;
        RECT 68.490 136.625 69.665 136.685 ;
        RECT 70.995 136.650 71.195 136.685 ;
        RECT 68.485 136.245 68.975 136.445 ;
        RECT 69.165 136.245 69.640 136.455 ;
        RECT 66.635 135.425 66.915 135.885 ;
        RECT 67.435 135.255 67.760 135.715 ;
        RECT 67.930 135.425 68.315 135.995 ;
        RECT 68.490 135.255 68.945 136.020 ;
        RECT 69.420 135.845 69.640 136.245 ;
        RECT 69.885 136.245 70.215 136.455 ;
        RECT 69.885 135.845 70.095 136.245 ;
        RECT 70.385 136.210 70.795 136.515 ;
        RECT 71.025 136.075 71.195 136.650 ;
        RECT 70.925 135.955 71.195 136.075 ;
        RECT 70.350 135.910 71.195 135.955 ;
        RECT 70.350 135.785 71.105 135.910 ;
        RECT 70.350 135.635 70.520 135.785 ;
        RECT 71.365 135.755 71.535 136.955 ;
        RECT 72.165 136.715 75.675 137.805 ;
        RECT 72.165 136.195 73.855 136.715 ;
        RECT 75.845 136.640 76.135 137.805 ;
        RECT 77.225 136.665 77.495 137.635 ;
        RECT 77.705 137.005 77.985 137.805 ;
        RECT 78.155 137.295 79.810 137.585 ;
        RECT 78.220 136.955 79.810 137.125 ;
        RECT 78.220 136.835 78.390 136.955 ;
        RECT 77.665 136.665 78.390 136.835 ;
        RECT 74.025 136.025 75.675 136.545 ;
        RECT 69.220 135.425 70.520 135.635 ;
        RECT 70.775 135.255 71.105 135.615 ;
        RECT 71.275 135.425 71.535 135.755 ;
        RECT 72.165 135.255 75.675 136.025 ;
        RECT 75.845 135.255 76.135 135.980 ;
        RECT 77.225 135.930 77.395 136.665 ;
        RECT 77.665 136.495 77.835 136.665 ;
        RECT 77.565 136.165 77.835 136.495 ;
        RECT 78.005 136.165 78.410 136.495 ;
        RECT 78.580 136.165 79.290 136.785 ;
        RECT 79.490 136.665 79.810 136.955 ;
        RECT 79.985 136.665 80.325 137.635 ;
        RECT 80.495 136.665 80.665 137.805 ;
        RECT 80.935 137.005 81.185 137.805 ;
        RECT 81.830 136.835 82.160 137.635 ;
        RECT 82.460 137.005 82.790 137.805 ;
        RECT 82.960 136.835 83.290 137.635 ;
        RECT 84.040 137.465 84.295 137.495 ;
        RECT 83.955 137.295 84.295 137.465 ;
        RECT 80.855 136.665 83.290 136.835 ;
        RECT 84.040 136.825 84.295 137.295 ;
        RECT 84.475 137.005 84.760 137.805 ;
        RECT 84.940 137.085 85.270 137.595 ;
        RECT 77.665 135.995 77.835 136.165 ;
        RECT 77.225 135.585 77.495 135.930 ;
        RECT 77.665 135.825 79.275 135.995 ;
        RECT 79.460 135.925 79.810 136.495 ;
        RECT 79.985 136.055 80.160 136.665 ;
        RECT 80.855 136.415 81.025 136.665 ;
        RECT 80.330 136.245 81.025 136.415 ;
        RECT 81.200 136.245 81.620 136.445 ;
        RECT 81.790 136.245 82.120 136.445 ;
        RECT 82.290 136.245 82.620 136.445 ;
        RECT 77.685 135.255 78.065 135.655 ;
        RECT 78.235 135.475 78.405 135.825 ;
        RECT 78.575 135.255 78.905 135.655 ;
        RECT 79.105 135.475 79.275 135.825 ;
        RECT 79.475 135.255 79.805 135.755 ;
        RECT 79.985 135.425 80.325 136.055 ;
        RECT 80.495 135.255 80.745 136.055 ;
        RECT 80.935 135.905 82.160 136.075 ;
        RECT 80.935 135.425 81.265 135.905 ;
        RECT 81.435 135.255 81.660 135.715 ;
        RECT 81.830 135.425 82.160 135.905 ;
        RECT 82.790 136.035 82.960 136.665 ;
        RECT 83.145 136.245 83.495 136.495 ;
        RECT 82.790 135.425 83.290 136.035 ;
        RECT 84.040 135.965 84.220 136.825 ;
        RECT 84.940 136.495 85.190 137.085 ;
        RECT 85.540 136.935 85.710 137.545 ;
        RECT 85.880 137.115 86.210 137.805 ;
        RECT 86.440 137.255 86.680 137.545 ;
        RECT 86.880 137.425 87.300 137.805 ;
        RECT 87.480 137.335 88.110 137.585 ;
        RECT 88.580 137.425 88.910 137.805 ;
        RECT 87.480 137.255 87.650 137.335 ;
        RECT 89.080 137.255 89.250 137.545 ;
        RECT 89.430 137.425 89.810 137.805 ;
        RECT 90.050 137.420 90.880 137.590 ;
        RECT 86.440 137.085 87.650 137.255 ;
        RECT 84.390 136.165 85.190 136.495 ;
        RECT 84.040 135.435 84.295 135.965 ;
        RECT 84.475 135.255 84.760 135.715 ;
        RECT 84.940 135.515 85.190 136.165 ;
        RECT 85.390 136.915 85.710 136.935 ;
        RECT 85.390 136.745 87.310 136.915 ;
        RECT 85.390 135.850 85.580 136.745 ;
        RECT 87.480 136.575 87.650 137.085 ;
        RECT 87.820 136.825 88.340 137.135 ;
        RECT 85.750 136.405 87.650 136.575 ;
        RECT 85.750 136.345 86.080 136.405 ;
        RECT 86.230 136.175 86.560 136.235 ;
        RECT 85.900 135.905 86.560 136.175 ;
        RECT 85.390 135.520 85.710 135.850 ;
        RECT 85.890 135.255 86.550 135.735 ;
        RECT 86.750 135.645 86.920 136.405 ;
        RECT 87.820 136.235 88.000 136.645 ;
        RECT 87.090 136.065 87.420 136.185 ;
        RECT 88.170 136.065 88.340 136.825 ;
        RECT 87.090 135.895 88.340 136.065 ;
        RECT 88.510 137.005 89.880 137.255 ;
        RECT 88.510 136.235 88.700 137.005 ;
        RECT 89.630 136.745 89.880 137.005 ;
        RECT 88.870 136.575 89.120 136.735 ;
        RECT 90.050 136.575 90.220 137.420 ;
        RECT 91.115 137.135 91.285 137.635 ;
        RECT 91.455 137.305 91.785 137.805 ;
        RECT 90.390 136.745 90.890 137.125 ;
        RECT 91.115 136.965 91.810 137.135 ;
        RECT 88.870 136.405 90.220 136.575 ;
        RECT 89.800 136.365 90.220 136.405 ;
        RECT 88.510 135.895 88.930 136.235 ;
        RECT 89.220 135.905 89.630 136.235 ;
        RECT 86.750 135.475 87.600 135.645 ;
        RECT 88.160 135.255 88.480 135.715 ;
        RECT 88.680 135.465 88.930 135.895 ;
        RECT 89.220 135.255 89.630 135.695 ;
        RECT 89.800 135.635 89.970 136.365 ;
        RECT 90.140 135.815 90.490 136.185 ;
        RECT 90.670 135.875 90.890 136.745 ;
        RECT 91.060 136.175 91.470 136.795 ;
        RECT 91.640 135.995 91.810 136.965 ;
        RECT 91.115 135.805 91.810 135.995 ;
        RECT 89.800 135.435 90.815 135.635 ;
        RECT 91.115 135.475 91.285 135.805 ;
        RECT 91.455 135.255 91.785 135.635 ;
        RECT 92.000 135.515 92.225 137.635 ;
        RECT 92.395 137.305 92.725 137.805 ;
        RECT 92.895 137.135 93.065 137.635 ;
        RECT 92.400 136.965 93.065 137.135 ;
        RECT 92.400 135.975 92.630 136.965 ;
        RECT 92.800 136.145 93.150 136.795 ;
        RECT 93.330 136.665 93.665 137.635 ;
        RECT 93.835 136.665 94.005 137.805 ;
        RECT 94.175 137.465 96.205 137.635 ;
        RECT 93.330 135.995 93.500 136.665 ;
        RECT 94.175 136.495 94.345 137.465 ;
        RECT 93.670 136.165 93.925 136.495 ;
        RECT 94.150 136.165 94.345 136.495 ;
        RECT 94.515 137.125 95.640 137.295 ;
        RECT 93.755 135.995 93.925 136.165 ;
        RECT 94.515 135.995 94.685 137.125 ;
        RECT 92.400 135.805 93.065 135.975 ;
        RECT 92.395 135.255 92.725 135.635 ;
        RECT 92.895 135.515 93.065 135.805 ;
        RECT 93.330 135.425 93.585 135.995 ;
        RECT 93.755 135.825 94.685 135.995 ;
        RECT 94.855 136.785 95.865 136.955 ;
        RECT 94.855 135.985 95.025 136.785 ;
        RECT 94.510 135.790 94.685 135.825 ;
        RECT 93.755 135.255 94.085 135.655 ;
        RECT 94.510 135.425 95.040 135.790 ;
        RECT 95.230 135.765 95.505 136.585 ;
        RECT 95.225 135.595 95.505 135.765 ;
        RECT 95.230 135.425 95.505 135.595 ;
        RECT 95.675 135.425 95.865 136.785 ;
        RECT 96.035 136.800 96.205 137.465 ;
        RECT 96.375 137.045 96.545 137.805 ;
        RECT 96.780 137.045 97.295 137.455 ;
        RECT 96.035 136.610 96.785 136.800 ;
        RECT 96.955 136.235 97.295 137.045 ;
        RECT 98.130 136.835 98.460 137.635 ;
        RECT 98.630 137.005 98.960 137.805 ;
        RECT 99.260 136.835 99.590 137.635 ;
        RECT 100.235 137.005 100.485 137.805 ;
        RECT 98.130 136.665 100.565 136.835 ;
        RECT 100.755 136.665 100.925 137.805 ;
        RECT 101.095 136.665 101.435 137.635 ;
        RECT 97.925 136.245 98.275 136.495 ;
        RECT 96.065 136.065 97.295 136.235 ;
        RECT 96.045 135.255 96.555 135.790 ;
        RECT 96.775 135.460 97.020 136.065 ;
        RECT 98.460 136.035 98.630 136.665 ;
        RECT 98.800 136.245 99.130 136.445 ;
        RECT 99.300 136.245 99.630 136.445 ;
        RECT 99.800 136.245 100.220 136.445 ;
        RECT 100.395 136.415 100.565 136.665 ;
        RECT 100.395 136.245 101.090 136.415 ;
        RECT 98.130 135.425 98.630 136.035 ;
        RECT 99.260 135.905 100.485 136.075 ;
        RECT 101.260 136.055 101.435 136.665 ;
        RECT 101.605 136.640 101.895 137.805 ;
        RECT 102.985 137.045 103.500 137.455 ;
        RECT 103.735 137.045 103.905 137.805 ;
        RECT 104.075 137.465 106.105 137.635 ;
        RECT 102.985 136.235 103.325 137.045 ;
        RECT 104.075 136.800 104.245 137.465 ;
        RECT 104.640 137.125 105.765 137.295 ;
        RECT 103.495 136.610 104.245 136.800 ;
        RECT 104.415 136.785 105.425 136.955 ;
        RECT 102.985 136.065 104.215 136.235 ;
        RECT 99.260 135.425 99.590 135.905 ;
        RECT 99.760 135.255 99.985 135.715 ;
        RECT 100.155 135.425 100.485 135.905 ;
        RECT 100.675 135.255 100.925 136.055 ;
        RECT 101.095 135.425 101.435 136.055 ;
        RECT 101.605 135.255 101.895 135.980 ;
        RECT 103.260 135.460 103.505 136.065 ;
        RECT 103.725 135.255 104.235 135.790 ;
        RECT 104.415 135.425 104.605 136.785 ;
        RECT 104.775 136.445 105.050 136.585 ;
        RECT 104.775 136.275 105.055 136.445 ;
        RECT 104.775 135.425 105.050 136.275 ;
        RECT 105.255 135.985 105.425 136.785 ;
        RECT 105.595 135.995 105.765 137.125 ;
        RECT 105.935 136.495 106.105 137.465 ;
        RECT 106.275 136.665 106.445 137.805 ;
        RECT 106.615 136.665 106.950 137.635 ;
        RECT 105.935 136.165 106.130 136.495 ;
        RECT 106.355 136.165 106.610 136.495 ;
        RECT 106.355 135.995 106.525 136.165 ;
        RECT 106.780 135.995 106.950 136.665 ;
        RECT 105.595 135.825 106.525 135.995 ;
        RECT 105.595 135.790 105.770 135.825 ;
        RECT 105.240 135.425 105.770 135.790 ;
        RECT 106.195 135.255 106.525 135.655 ;
        RECT 106.695 135.425 106.950 135.995 ;
        RECT 107.125 136.730 107.395 137.635 ;
        RECT 107.565 137.045 107.895 137.805 ;
        RECT 108.075 136.875 108.245 137.635 ;
        RECT 107.125 135.930 107.295 136.730 ;
        RECT 107.580 136.705 108.245 136.875 ;
        RECT 109.425 137.045 109.940 137.455 ;
        RECT 110.175 137.045 110.345 137.805 ;
        RECT 110.515 137.465 112.545 137.635 ;
        RECT 107.580 136.560 107.750 136.705 ;
        RECT 107.465 136.230 107.750 136.560 ;
        RECT 107.580 135.975 107.750 136.230 ;
        RECT 107.985 136.155 108.315 136.525 ;
        RECT 109.425 136.235 109.765 137.045 ;
        RECT 110.515 136.800 110.685 137.465 ;
        RECT 111.080 137.125 112.205 137.295 ;
        RECT 109.935 136.610 110.685 136.800 ;
        RECT 110.855 136.785 111.865 136.955 ;
        RECT 109.425 136.065 110.655 136.235 ;
        RECT 107.125 135.425 107.385 135.930 ;
        RECT 107.580 135.805 108.245 135.975 ;
        RECT 107.565 135.255 107.895 135.635 ;
        RECT 108.075 135.425 108.245 135.805 ;
        RECT 109.700 135.460 109.945 136.065 ;
        RECT 110.165 135.255 110.675 135.790 ;
        RECT 110.855 135.425 111.045 136.785 ;
        RECT 111.215 136.445 111.490 136.585 ;
        RECT 111.215 136.275 111.495 136.445 ;
        RECT 111.215 135.425 111.490 136.275 ;
        RECT 111.695 135.985 111.865 136.785 ;
        RECT 112.035 135.995 112.205 137.125 ;
        RECT 112.375 136.495 112.545 137.465 ;
        RECT 112.715 136.665 112.885 137.805 ;
        RECT 113.055 136.665 113.390 137.635 ;
        RECT 112.375 136.165 112.570 136.495 ;
        RECT 112.795 136.165 113.050 136.495 ;
        RECT 112.795 135.995 112.965 136.165 ;
        RECT 113.220 135.995 113.390 136.665 ;
        RECT 113.940 136.825 114.195 137.495 ;
        RECT 114.375 137.005 114.660 137.805 ;
        RECT 114.840 137.085 115.170 137.595 ;
        RECT 113.940 136.105 114.120 136.825 ;
        RECT 114.840 136.495 115.090 137.085 ;
        RECT 115.440 136.935 115.610 137.545 ;
        RECT 115.780 137.115 116.110 137.805 ;
        RECT 116.340 137.255 116.580 137.545 ;
        RECT 116.780 137.425 117.200 137.805 ;
        RECT 117.380 137.335 118.010 137.585 ;
        RECT 118.480 137.425 118.810 137.805 ;
        RECT 117.380 137.255 117.550 137.335 ;
        RECT 118.980 137.255 119.150 137.545 ;
        RECT 119.330 137.425 119.710 137.805 ;
        RECT 119.950 137.420 120.780 137.590 ;
        RECT 116.340 137.085 117.550 137.255 ;
        RECT 114.290 136.165 115.090 136.495 ;
        RECT 112.035 135.825 112.965 135.995 ;
        RECT 112.035 135.790 112.210 135.825 ;
        RECT 111.680 135.425 112.210 135.790 ;
        RECT 112.635 135.255 112.965 135.655 ;
        RECT 113.135 135.425 113.390 135.995 ;
        RECT 113.855 135.965 114.120 136.105 ;
        RECT 113.855 135.935 114.195 135.965 ;
        RECT 113.940 135.435 114.195 135.935 ;
        RECT 114.375 135.255 114.660 135.715 ;
        RECT 114.840 135.515 115.090 136.165 ;
        RECT 115.290 136.915 115.610 136.935 ;
        RECT 115.290 136.745 117.210 136.915 ;
        RECT 115.290 135.850 115.480 136.745 ;
        RECT 117.380 136.575 117.550 137.085 ;
        RECT 117.720 136.825 118.240 137.135 ;
        RECT 115.650 136.405 117.550 136.575 ;
        RECT 115.650 136.345 115.980 136.405 ;
        RECT 116.130 136.175 116.460 136.235 ;
        RECT 115.800 135.905 116.460 136.175 ;
        RECT 115.290 135.520 115.610 135.850 ;
        RECT 115.790 135.255 116.450 135.735 ;
        RECT 116.650 135.645 116.820 136.405 ;
        RECT 117.720 136.235 117.900 136.645 ;
        RECT 116.990 136.065 117.320 136.185 ;
        RECT 118.070 136.065 118.240 136.825 ;
        RECT 116.990 135.895 118.240 136.065 ;
        RECT 118.410 137.005 119.780 137.255 ;
        RECT 118.410 136.235 118.600 137.005 ;
        RECT 119.530 136.745 119.780 137.005 ;
        RECT 118.770 136.575 119.020 136.735 ;
        RECT 119.950 136.575 120.120 137.420 ;
        RECT 121.015 137.135 121.185 137.635 ;
        RECT 121.355 137.305 121.685 137.805 ;
        RECT 120.290 136.745 120.790 137.125 ;
        RECT 121.015 136.965 121.710 137.135 ;
        RECT 118.770 136.405 120.120 136.575 ;
        RECT 119.700 136.365 120.120 136.405 ;
        RECT 118.410 135.895 118.830 136.235 ;
        RECT 119.120 135.905 119.530 136.235 ;
        RECT 116.650 135.475 117.500 135.645 ;
        RECT 118.060 135.255 118.380 135.715 ;
        RECT 118.580 135.465 118.830 135.895 ;
        RECT 119.120 135.255 119.530 135.695 ;
        RECT 119.700 135.635 119.870 136.365 ;
        RECT 120.040 135.815 120.390 136.185 ;
        RECT 120.570 135.875 120.790 136.745 ;
        RECT 120.960 136.175 121.370 136.795 ;
        RECT 121.540 135.995 121.710 136.965 ;
        RECT 121.015 135.805 121.710 135.995 ;
        RECT 119.700 135.435 120.715 135.635 ;
        RECT 121.015 135.475 121.185 135.805 ;
        RECT 121.355 135.255 121.685 135.635 ;
        RECT 121.900 135.515 122.125 137.635 ;
        RECT 122.295 137.305 122.625 137.805 ;
        RECT 122.795 137.135 122.965 137.635 ;
        RECT 122.300 136.965 122.965 137.135 ;
        RECT 122.300 135.975 122.530 136.965 ;
        RECT 123.315 136.875 123.485 137.635 ;
        RECT 123.665 137.045 123.995 137.805 ;
        RECT 122.700 136.145 123.050 136.795 ;
        RECT 123.315 136.705 123.980 136.875 ;
        RECT 124.165 136.730 124.435 137.635 ;
        RECT 123.810 136.560 123.980 136.705 ;
        RECT 123.245 136.155 123.575 136.525 ;
        RECT 123.810 136.230 124.095 136.560 ;
        RECT 123.810 135.975 123.980 136.230 ;
        RECT 122.300 135.805 122.965 135.975 ;
        RECT 122.295 135.255 122.625 135.635 ;
        RECT 122.795 135.515 122.965 135.805 ;
        RECT 123.315 135.805 123.980 135.975 ;
        RECT 124.265 135.930 124.435 136.730 ;
        RECT 124.605 136.715 126.275 137.805 ;
        RECT 126.445 136.715 127.655 137.805 ;
        RECT 124.605 136.195 125.355 136.715 ;
        RECT 125.525 136.025 126.275 136.545 ;
        RECT 126.445 136.175 126.965 136.715 ;
        RECT 123.315 135.425 123.485 135.805 ;
        RECT 123.665 135.255 123.995 135.635 ;
        RECT 124.175 135.425 124.435 135.930 ;
        RECT 124.605 135.255 126.275 136.025 ;
        RECT 127.135 136.005 127.655 136.545 ;
        RECT 126.445 135.255 127.655 136.005 ;
        RECT 14.580 135.085 127.740 135.255 ;
        RECT 14.665 134.335 15.875 135.085 ;
        RECT 14.665 133.795 15.185 134.335 ;
        RECT 16.565 134.265 16.775 135.085 ;
        RECT 16.945 134.285 17.275 134.915 ;
        RECT 15.355 133.625 15.875 134.165 ;
        RECT 16.945 133.685 17.195 134.285 ;
        RECT 17.445 134.265 17.675 135.085 ;
        RECT 17.975 134.535 18.145 134.915 ;
        RECT 18.325 134.705 18.655 135.085 ;
        RECT 17.975 134.365 18.640 134.535 ;
        RECT 18.835 134.410 19.095 134.915 ;
        RECT 17.365 133.845 17.695 134.095 ;
        RECT 17.905 133.815 18.235 134.185 ;
        RECT 18.470 134.110 18.640 134.365 ;
        RECT 18.470 133.780 18.755 134.110 ;
        RECT 14.665 132.535 15.875 133.625 ;
        RECT 16.565 132.535 16.775 133.675 ;
        RECT 16.945 132.705 17.275 133.685 ;
        RECT 17.445 132.535 17.675 133.675 ;
        RECT 18.470 133.635 18.640 133.780 ;
        RECT 17.975 133.465 18.640 133.635 ;
        RECT 18.925 133.610 19.095 134.410 ;
        RECT 19.305 134.265 19.535 135.085 ;
        RECT 19.705 134.285 20.035 134.915 ;
        RECT 19.285 133.845 19.615 134.095 ;
        RECT 19.785 133.685 20.035 134.285 ;
        RECT 20.205 134.265 20.415 135.085 ;
        RECT 21.020 134.745 21.275 134.905 ;
        RECT 20.935 134.575 21.275 134.745 ;
        RECT 21.455 134.625 21.740 135.085 ;
        RECT 21.020 134.375 21.275 134.575 ;
        RECT 17.975 132.705 18.145 133.465 ;
        RECT 18.325 132.535 18.655 133.295 ;
        RECT 18.825 132.705 19.095 133.610 ;
        RECT 19.305 132.535 19.535 133.675 ;
        RECT 19.705 132.705 20.035 133.685 ;
        RECT 20.205 132.535 20.415 133.675 ;
        RECT 21.020 133.515 21.200 134.375 ;
        RECT 21.920 134.175 22.170 134.825 ;
        RECT 21.370 133.845 22.170 134.175 ;
        RECT 21.020 132.845 21.275 133.515 ;
        RECT 21.455 132.535 21.740 133.335 ;
        RECT 21.920 133.255 22.170 133.845 ;
        RECT 22.370 134.490 22.690 134.820 ;
        RECT 22.870 134.605 23.530 135.085 ;
        RECT 23.730 134.695 24.580 134.865 ;
        RECT 22.370 133.595 22.560 134.490 ;
        RECT 22.880 134.165 23.540 134.435 ;
        RECT 23.210 134.105 23.540 134.165 ;
        RECT 22.730 133.935 23.060 133.995 ;
        RECT 23.730 133.935 23.900 134.695 ;
        RECT 25.140 134.625 25.460 135.085 ;
        RECT 25.660 134.445 25.910 134.875 ;
        RECT 26.200 134.645 26.610 135.085 ;
        RECT 26.780 134.705 27.795 134.905 ;
        RECT 24.070 134.275 25.320 134.445 ;
        RECT 24.070 134.155 24.400 134.275 ;
        RECT 22.730 133.765 24.630 133.935 ;
        RECT 22.370 133.425 24.290 133.595 ;
        RECT 22.370 133.405 22.690 133.425 ;
        RECT 21.920 132.745 22.250 133.255 ;
        RECT 22.520 132.795 22.690 133.405 ;
        RECT 24.460 133.255 24.630 133.765 ;
        RECT 24.800 133.695 24.980 134.105 ;
        RECT 25.150 133.515 25.320 134.275 ;
        RECT 22.860 132.535 23.190 133.225 ;
        RECT 23.420 133.085 24.630 133.255 ;
        RECT 24.800 133.205 25.320 133.515 ;
        RECT 25.490 134.105 25.910 134.445 ;
        RECT 26.200 134.105 26.610 134.435 ;
        RECT 25.490 133.335 25.680 134.105 ;
        RECT 26.780 133.975 26.950 134.705 ;
        RECT 28.095 134.535 28.265 134.865 ;
        RECT 28.435 134.705 28.765 135.085 ;
        RECT 27.120 134.155 27.470 134.525 ;
        RECT 26.780 133.935 27.200 133.975 ;
        RECT 25.850 133.765 27.200 133.935 ;
        RECT 25.850 133.605 26.100 133.765 ;
        RECT 26.610 133.335 26.860 133.595 ;
        RECT 25.490 133.085 26.860 133.335 ;
        RECT 23.420 132.795 23.660 133.085 ;
        RECT 24.460 133.005 24.630 133.085 ;
        RECT 23.860 132.535 24.280 132.915 ;
        RECT 24.460 132.755 25.090 133.005 ;
        RECT 25.560 132.535 25.890 132.915 ;
        RECT 26.060 132.795 26.230 133.085 ;
        RECT 27.030 132.920 27.200 133.765 ;
        RECT 27.650 133.595 27.870 134.465 ;
        RECT 28.095 134.345 28.790 134.535 ;
        RECT 27.370 133.215 27.870 133.595 ;
        RECT 28.040 133.545 28.450 134.165 ;
        RECT 28.620 133.375 28.790 134.345 ;
        RECT 28.095 133.205 28.790 133.375 ;
        RECT 26.410 132.535 26.790 132.915 ;
        RECT 27.030 132.750 27.860 132.920 ;
        RECT 28.095 132.705 28.265 133.205 ;
        RECT 28.435 132.535 28.765 133.035 ;
        RECT 28.980 132.705 29.205 134.825 ;
        RECT 29.375 134.705 29.705 135.085 ;
        RECT 29.875 134.535 30.045 134.825 ;
        RECT 29.380 134.365 30.045 134.535 ;
        RECT 30.965 134.455 31.295 134.815 ;
        RECT 31.915 134.625 32.165 135.085 ;
        RECT 32.335 134.625 32.895 134.915 ;
        RECT 29.380 133.375 29.610 134.365 ;
        RECT 30.965 134.265 32.355 134.455 ;
        RECT 29.780 133.545 30.130 134.195 ;
        RECT 32.185 134.175 32.355 134.265 ;
        RECT 30.780 133.845 31.455 134.095 ;
        RECT 31.675 133.845 32.015 134.095 ;
        RECT 32.185 133.845 32.475 134.175 ;
        RECT 30.780 133.485 31.045 133.845 ;
        RECT 32.185 133.595 32.355 133.845 ;
        RECT 31.415 133.425 32.355 133.595 ;
        RECT 29.380 133.205 30.045 133.375 ;
        RECT 29.375 132.535 29.705 133.035 ;
        RECT 29.875 132.705 30.045 133.205 ;
        RECT 30.965 132.535 31.245 133.205 ;
        RECT 31.415 132.875 31.715 133.425 ;
        RECT 32.645 133.255 32.895 134.625 ;
        RECT 33.340 134.275 33.585 134.880 ;
        RECT 33.805 134.550 34.315 135.085 ;
        RECT 31.915 132.535 32.245 133.255 ;
        RECT 32.435 132.705 32.895 133.255 ;
        RECT 33.065 134.105 34.295 134.275 ;
        RECT 33.065 133.295 33.405 134.105 ;
        RECT 33.575 133.540 34.325 133.730 ;
        RECT 33.065 132.885 33.580 133.295 ;
        RECT 33.815 132.535 33.985 133.295 ;
        RECT 34.155 132.875 34.325 133.540 ;
        RECT 34.495 133.555 34.685 134.915 ;
        RECT 34.855 134.065 35.130 134.915 ;
        RECT 35.320 134.550 35.850 134.915 ;
        RECT 36.275 134.685 36.605 135.085 ;
        RECT 35.675 134.515 35.850 134.550 ;
        RECT 34.855 133.895 35.135 134.065 ;
        RECT 34.855 133.755 35.130 133.895 ;
        RECT 35.335 133.555 35.505 134.355 ;
        RECT 34.495 133.385 35.505 133.555 ;
        RECT 35.675 134.345 36.605 134.515 ;
        RECT 36.775 134.345 37.030 134.915 ;
        RECT 37.205 134.360 37.495 135.085 ;
        RECT 35.675 133.215 35.845 134.345 ;
        RECT 36.435 134.175 36.605 134.345 ;
        RECT 34.720 133.045 35.845 133.215 ;
        RECT 36.015 133.845 36.210 134.175 ;
        RECT 36.435 133.845 36.690 134.175 ;
        RECT 36.015 132.875 36.185 133.845 ;
        RECT 36.860 133.675 37.030 134.345 ;
        RECT 37.665 134.315 39.335 135.085 ;
        RECT 39.515 134.585 39.845 135.085 ;
        RECT 40.045 134.515 40.215 134.865 ;
        RECT 40.415 134.685 40.745 135.085 ;
        RECT 40.915 134.515 41.085 134.865 ;
        RECT 41.255 134.685 41.635 135.085 ;
        RECT 34.155 132.705 36.185 132.875 ;
        RECT 36.355 132.535 36.525 133.675 ;
        RECT 36.695 132.705 37.030 133.675 ;
        RECT 37.205 132.535 37.495 133.700 ;
        RECT 37.665 133.625 38.415 134.145 ;
        RECT 38.585 133.795 39.335 134.315 ;
        RECT 39.510 133.845 39.860 134.415 ;
        RECT 40.045 134.345 41.655 134.515 ;
        RECT 41.825 134.410 42.095 134.755 ;
        RECT 42.275 134.585 42.605 135.085 ;
        RECT 42.805 134.515 42.975 134.865 ;
        RECT 43.175 134.685 43.505 135.085 ;
        RECT 43.675 134.515 43.845 134.865 ;
        RECT 44.015 134.685 44.395 135.085 ;
        RECT 41.485 134.175 41.655 134.345 ;
        RECT 37.665 132.535 39.335 133.625 ;
        RECT 39.510 133.385 39.830 133.675 ;
        RECT 40.030 133.555 40.740 134.175 ;
        RECT 40.910 133.845 41.315 134.175 ;
        RECT 41.485 133.845 41.755 134.175 ;
        RECT 41.485 133.675 41.655 133.845 ;
        RECT 41.925 133.675 42.095 134.410 ;
        RECT 42.270 133.845 42.620 134.415 ;
        RECT 42.805 134.345 44.415 134.515 ;
        RECT 44.585 134.410 44.855 134.755 ;
        RECT 44.245 134.175 44.415 134.345 ;
        RECT 40.930 133.505 41.655 133.675 ;
        RECT 40.930 133.385 41.100 133.505 ;
        RECT 39.510 133.215 41.100 133.385 ;
        RECT 39.510 132.755 41.165 133.045 ;
        RECT 41.335 132.535 41.615 133.335 ;
        RECT 41.825 132.705 42.095 133.675 ;
        RECT 42.270 133.385 42.590 133.675 ;
        RECT 42.790 133.555 43.500 134.175 ;
        RECT 43.670 133.845 44.075 134.175 ;
        RECT 44.245 133.845 44.515 134.175 ;
        RECT 44.245 133.675 44.415 133.845 ;
        RECT 44.685 133.675 44.855 134.410 ;
        RECT 43.690 133.505 44.415 133.675 ;
        RECT 43.690 133.385 43.860 133.505 ;
        RECT 42.270 133.215 43.860 133.385 ;
        RECT 42.270 132.755 43.925 133.045 ;
        RECT 44.095 132.535 44.375 133.335 ;
        RECT 44.585 132.705 44.855 133.675 ;
        RECT 45.025 134.285 45.365 134.915 ;
        RECT 45.535 134.285 45.785 135.085 ;
        RECT 45.975 134.435 46.305 134.915 ;
        RECT 46.475 134.625 46.700 135.085 ;
        RECT 46.870 134.435 47.200 134.915 ;
        RECT 45.025 133.725 45.200 134.285 ;
        RECT 45.975 134.265 47.200 134.435 ;
        RECT 47.830 134.305 48.330 134.915 ;
        RECT 45.370 133.925 46.065 134.095 ;
        RECT 45.025 133.675 45.255 133.725 ;
        RECT 45.895 133.675 46.065 133.925 ;
        RECT 46.240 133.895 46.660 134.095 ;
        RECT 46.830 133.895 47.160 134.095 ;
        RECT 47.330 133.895 47.660 134.095 ;
        RECT 47.830 133.675 48.000 134.305 ;
        RECT 48.705 134.285 49.045 134.915 ;
        RECT 49.215 134.285 49.465 135.085 ;
        RECT 49.655 134.435 49.985 134.915 ;
        RECT 50.155 134.625 50.380 135.085 ;
        RECT 50.550 134.435 50.880 134.915 ;
        RECT 48.705 134.235 48.935 134.285 ;
        RECT 49.655 134.265 50.880 134.435 ;
        RECT 51.510 134.305 52.010 134.915 ;
        RECT 52.760 134.745 53.015 134.905 ;
        RECT 52.675 134.575 53.015 134.745 ;
        RECT 53.195 134.625 53.480 135.085 ;
        RECT 52.760 134.375 53.015 134.575 ;
        RECT 48.185 133.845 48.535 134.095 ;
        RECT 48.705 133.675 48.880 134.235 ;
        RECT 49.050 133.925 49.745 134.095 ;
        RECT 49.575 133.675 49.745 133.925 ;
        RECT 49.920 133.895 50.340 134.095 ;
        RECT 50.510 133.895 50.840 134.095 ;
        RECT 51.010 133.895 51.340 134.095 ;
        RECT 51.510 133.675 51.680 134.305 ;
        RECT 51.865 133.845 52.215 134.095 ;
        RECT 45.025 132.705 45.365 133.675 ;
        RECT 45.535 132.535 45.705 133.675 ;
        RECT 45.895 133.505 48.330 133.675 ;
        RECT 45.975 132.535 46.225 133.335 ;
        RECT 46.870 132.705 47.200 133.505 ;
        RECT 47.500 132.535 47.830 133.335 ;
        RECT 48.000 132.705 48.330 133.505 ;
        RECT 48.705 132.705 49.045 133.675 ;
        RECT 49.215 132.535 49.385 133.675 ;
        RECT 49.575 133.505 52.010 133.675 ;
        RECT 49.655 132.535 49.905 133.335 ;
        RECT 50.550 132.705 50.880 133.505 ;
        RECT 51.180 132.535 51.510 133.335 ;
        RECT 51.680 132.705 52.010 133.505 ;
        RECT 52.760 133.515 52.940 134.375 ;
        RECT 53.660 134.175 53.910 134.825 ;
        RECT 53.110 133.845 53.910 134.175 ;
        RECT 52.760 132.845 53.015 133.515 ;
        RECT 53.195 132.535 53.480 133.335 ;
        RECT 53.660 133.255 53.910 133.845 ;
        RECT 54.110 134.490 54.430 134.820 ;
        RECT 54.610 134.605 55.270 135.085 ;
        RECT 55.470 134.695 56.320 134.865 ;
        RECT 54.110 133.595 54.300 134.490 ;
        RECT 54.620 134.165 55.280 134.435 ;
        RECT 54.950 134.105 55.280 134.165 ;
        RECT 54.470 133.935 54.800 133.995 ;
        RECT 55.470 133.935 55.640 134.695 ;
        RECT 56.880 134.625 57.200 135.085 ;
        RECT 57.400 134.445 57.650 134.875 ;
        RECT 57.940 134.645 58.350 135.085 ;
        RECT 58.520 134.705 59.535 134.905 ;
        RECT 55.810 134.275 57.060 134.445 ;
        RECT 55.810 134.155 56.140 134.275 ;
        RECT 54.470 133.765 56.370 133.935 ;
        RECT 54.110 133.425 56.030 133.595 ;
        RECT 54.110 133.405 54.430 133.425 ;
        RECT 53.660 132.745 53.990 133.255 ;
        RECT 54.260 132.795 54.430 133.405 ;
        RECT 56.200 133.255 56.370 133.765 ;
        RECT 56.540 133.695 56.720 134.105 ;
        RECT 56.890 133.515 57.060 134.275 ;
        RECT 54.600 132.535 54.930 133.225 ;
        RECT 55.160 133.085 56.370 133.255 ;
        RECT 56.540 133.205 57.060 133.515 ;
        RECT 57.230 134.105 57.650 134.445 ;
        RECT 57.940 134.105 58.350 134.435 ;
        RECT 57.230 133.335 57.420 134.105 ;
        RECT 58.520 133.975 58.690 134.705 ;
        RECT 59.835 134.535 60.005 134.865 ;
        RECT 60.175 134.705 60.505 135.085 ;
        RECT 58.860 134.155 59.210 134.525 ;
        RECT 58.520 133.935 58.940 133.975 ;
        RECT 57.590 133.765 58.940 133.935 ;
        RECT 57.590 133.605 57.840 133.765 ;
        RECT 58.350 133.335 58.600 133.595 ;
        RECT 57.230 133.085 58.600 133.335 ;
        RECT 55.160 132.795 55.400 133.085 ;
        RECT 56.200 133.005 56.370 133.085 ;
        RECT 55.600 132.535 56.020 132.915 ;
        RECT 56.200 132.755 56.830 133.005 ;
        RECT 57.300 132.535 57.630 132.915 ;
        RECT 57.800 132.795 57.970 133.085 ;
        RECT 58.770 132.920 58.940 133.765 ;
        RECT 59.390 133.595 59.610 134.465 ;
        RECT 59.835 134.345 60.530 134.535 ;
        RECT 59.110 133.215 59.610 133.595 ;
        RECT 59.780 133.545 60.190 134.165 ;
        RECT 60.360 133.375 60.530 134.345 ;
        RECT 59.835 133.205 60.530 133.375 ;
        RECT 58.150 132.535 58.530 132.915 ;
        RECT 58.770 132.750 59.600 132.920 ;
        RECT 59.835 132.705 60.005 133.205 ;
        RECT 60.175 132.535 60.505 133.035 ;
        RECT 60.720 132.705 60.945 134.825 ;
        RECT 61.115 134.705 61.445 135.085 ;
        RECT 61.615 134.535 61.785 134.825 ;
        RECT 61.120 134.365 61.785 134.535 ;
        RECT 61.120 133.375 61.350 134.365 ;
        RECT 62.965 134.360 63.255 135.085 ;
        RECT 63.425 134.285 63.765 134.915 ;
        RECT 63.935 134.285 64.185 135.085 ;
        RECT 64.375 134.435 64.705 134.915 ;
        RECT 64.875 134.625 65.100 135.085 ;
        RECT 65.270 134.435 65.600 134.915 ;
        RECT 61.520 133.545 61.870 134.195 ;
        RECT 63.425 133.725 63.600 134.285 ;
        RECT 64.375 134.265 65.600 134.435 ;
        RECT 66.230 134.305 66.730 134.915 ;
        RECT 68.030 134.540 73.375 135.085 ;
        RECT 73.550 134.540 78.895 135.085 ;
        RECT 79.075 134.585 79.405 135.085 ;
        RECT 63.770 133.925 64.465 134.095 ;
        RECT 61.120 133.205 61.785 133.375 ;
        RECT 61.115 132.535 61.445 133.035 ;
        RECT 61.615 132.705 61.785 133.205 ;
        RECT 62.965 132.535 63.255 133.700 ;
        RECT 63.425 133.675 63.655 133.725 ;
        RECT 64.295 133.675 64.465 133.925 ;
        RECT 64.640 133.895 65.060 134.095 ;
        RECT 65.230 133.895 65.560 134.095 ;
        RECT 65.730 133.895 66.060 134.095 ;
        RECT 66.230 133.675 66.400 134.305 ;
        RECT 66.585 133.845 66.935 134.095 ;
        RECT 63.425 132.705 63.765 133.675 ;
        RECT 63.935 132.535 64.105 133.675 ;
        RECT 64.295 133.505 66.730 133.675 ;
        RECT 64.375 132.535 64.625 133.335 ;
        RECT 65.270 132.705 65.600 133.505 ;
        RECT 65.900 132.535 66.230 133.335 ;
        RECT 66.400 132.705 66.730 133.505 ;
        RECT 69.620 132.970 69.970 134.220 ;
        RECT 71.450 133.710 71.790 134.540 ;
        RECT 75.140 132.970 75.490 134.220 ;
        RECT 76.970 133.710 77.310 134.540 ;
        RECT 79.605 134.515 79.775 134.865 ;
        RECT 79.975 134.685 80.305 135.085 ;
        RECT 80.475 134.515 80.645 134.865 ;
        RECT 80.815 134.685 81.195 135.085 ;
        RECT 79.070 133.845 79.420 134.415 ;
        RECT 79.605 134.345 81.215 134.515 ;
        RECT 81.385 134.410 81.655 134.755 ;
        RECT 81.830 134.540 87.175 135.085 ;
        RECT 81.045 134.175 81.215 134.345 ;
        RECT 79.070 133.385 79.390 133.675 ;
        RECT 79.590 133.555 80.300 134.175 ;
        RECT 80.470 133.845 80.875 134.175 ;
        RECT 81.045 133.845 81.315 134.175 ;
        RECT 81.045 133.675 81.215 133.845 ;
        RECT 81.485 133.675 81.655 134.410 ;
        RECT 80.490 133.505 81.215 133.675 ;
        RECT 80.490 133.385 80.660 133.505 ;
        RECT 79.070 133.215 80.660 133.385 ;
        RECT 68.030 132.535 73.375 132.970 ;
        RECT 73.550 132.535 78.895 132.970 ;
        RECT 79.070 132.755 80.725 133.045 ;
        RECT 80.895 132.535 81.175 133.335 ;
        RECT 81.385 132.705 81.655 133.675 ;
        RECT 83.420 132.970 83.770 134.220 ;
        RECT 85.250 133.710 85.590 134.540 ;
        RECT 87.405 134.265 87.615 135.085 ;
        RECT 87.785 134.285 88.115 134.915 ;
        RECT 87.785 133.685 88.035 134.285 ;
        RECT 88.285 134.265 88.515 135.085 ;
        RECT 88.725 134.360 89.015 135.085 ;
        RECT 89.560 134.375 89.815 134.905 ;
        RECT 89.995 134.625 90.280 135.085 ;
        RECT 88.205 133.845 88.535 134.095 ;
        RECT 89.560 133.725 89.740 134.375 ;
        RECT 90.460 134.175 90.710 134.825 ;
        RECT 89.910 133.845 90.710 134.175 ;
        RECT 81.830 132.535 87.175 132.970 ;
        RECT 87.405 132.535 87.615 133.675 ;
        RECT 87.785 132.705 88.115 133.685 ;
        RECT 88.285 132.535 88.515 133.675 ;
        RECT 88.725 132.535 89.015 133.700 ;
        RECT 89.475 133.555 89.740 133.725 ;
        RECT 89.560 133.515 89.740 133.555 ;
        RECT 89.560 132.845 89.815 133.515 ;
        RECT 89.995 132.535 90.280 133.335 ;
        RECT 90.460 133.255 90.710 133.845 ;
        RECT 90.910 134.490 91.230 134.820 ;
        RECT 91.410 134.605 92.070 135.085 ;
        RECT 92.270 134.695 93.120 134.865 ;
        RECT 90.910 133.595 91.100 134.490 ;
        RECT 91.420 134.165 92.080 134.435 ;
        RECT 91.750 134.105 92.080 134.165 ;
        RECT 91.270 133.935 91.600 133.995 ;
        RECT 92.270 133.935 92.440 134.695 ;
        RECT 93.680 134.625 94.000 135.085 ;
        RECT 94.200 134.445 94.450 134.875 ;
        RECT 94.740 134.645 95.150 135.085 ;
        RECT 95.320 134.705 96.335 134.905 ;
        RECT 92.610 134.275 93.860 134.445 ;
        RECT 92.610 134.155 92.940 134.275 ;
        RECT 91.270 133.765 93.170 133.935 ;
        RECT 90.910 133.425 92.830 133.595 ;
        RECT 90.910 133.405 91.230 133.425 ;
        RECT 90.460 132.745 90.790 133.255 ;
        RECT 91.060 132.795 91.230 133.405 ;
        RECT 93.000 133.255 93.170 133.765 ;
        RECT 93.340 133.695 93.520 134.105 ;
        RECT 93.690 133.515 93.860 134.275 ;
        RECT 91.400 132.535 91.730 133.225 ;
        RECT 91.960 133.085 93.170 133.255 ;
        RECT 93.340 133.205 93.860 133.515 ;
        RECT 94.030 134.105 94.450 134.445 ;
        RECT 94.740 134.105 95.150 134.435 ;
        RECT 94.030 133.335 94.220 134.105 ;
        RECT 95.320 133.975 95.490 134.705 ;
        RECT 96.635 134.535 96.805 134.865 ;
        RECT 96.975 134.705 97.305 135.085 ;
        RECT 95.660 134.155 96.010 134.525 ;
        RECT 95.320 133.935 95.740 133.975 ;
        RECT 94.390 133.765 95.740 133.935 ;
        RECT 94.390 133.605 94.640 133.765 ;
        RECT 95.150 133.335 95.400 133.595 ;
        RECT 94.030 133.085 95.400 133.335 ;
        RECT 91.960 132.795 92.200 133.085 ;
        RECT 93.000 133.005 93.170 133.085 ;
        RECT 92.400 132.535 92.820 132.915 ;
        RECT 93.000 132.755 93.630 133.005 ;
        RECT 94.100 132.535 94.430 132.915 ;
        RECT 94.600 132.795 94.770 133.085 ;
        RECT 95.570 132.920 95.740 133.765 ;
        RECT 96.190 133.595 96.410 134.465 ;
        RECT 96.635 134.345 97.330 134.535 ;
        RECT 95.910 133.215 96.410 133.595 ;
        RECT 96.580 133.545 96.990 134.165 ;
        RECT 97.160 133.375 97.330 134.345 ;
        RECT 96.635 133.205 97.330 133.375 ;
        RECT 94.950 132.535 95.330 132.915 ;
        RECT 95.570 132.750 96.400 132.920 ;
        RECT 96.635 132.705 96.805 133.205 ;
        RECT 96.975 132.535 97.305 133.035 ;
        RECT 97.520 132.705 97.745 134.825 ;
        RECT 97.915 134.705 98.245 135.085 ;
        RECT 98.415 134.535 98.585 134.825 ;
        RECT 97.920 134.365 98.585 134.535 ;
        RECT 98.845 134.410 99.115 134.755 ;
        RECT 99.305 134.685 99.685 135.085 ;
        RECT 99.855 134.515 100.025 134.865 ;
        RECT 100.195 134.685 100.525 135.085 ;
        RECT 100.725 134.515 100.895 134.865 ;
        RECT 101.095 134.585 101.425 135.085 ;
        RECT 97.920 133.375 98.150 134.365 ;
        RECT 98.320 133.545 98.670 134.195 ;
        RECT 98.845 133.675 99.015 134.410 ;
        RECT 99.285 134.345 100.895 134.515 ;
        RECT 99.285 134.175 99.455 134.345 ;
        RECT 99.185 133.845 99.455 134.175 ;
        RECT 99.625 133.845 100.030 134.175 ;
        RECT 99.285 133.675 99.455 133.845 ;
        RECT 100.200 133.725 100.910 134.175 ;
        RECT 101.080 133.845 101.430 134.415 ;
        RECT 101.665 134.265 101.875 135.085 ;
        RECT 102.045 134.285 102.375 134.915 ;
        RECT 97.920 133.205 98.585 133.375 ;
        RECT 97.915 132.535 98.245 133.035 ;
        RECT 98.415 132.705 98.585 133.205 ;
        RECT 98.845 132.705 99.115 133.675 ;
        RECT 99.285 133.505 100.010 133.675 ;
        RECT 100.200 133.555 100.915 133.725 ;
        RECT 102.045 133.685 102.295 134.285 ;
        RECT 102.545 134.265 102.775 135.085 ;
        RECT 103.445 134.410 103.715 134.755 ;
        RECT 103.905 134.685 104.285 135.085 ;
        RECT 104.455 134.515 104.625 134.865 ;
        RECT 104.795 134.685 105.125 135.085 ;
        RECT 105.325 134.515 105.495 134.865 ;
        RECT 105.695 134.585 106.025 135.085 ;
        RECT 102.465 133.845 102.795 134.095 ;
        RECT 99.840 133.385 100.010 133.505 ;
        RECT 101.110 133.385 101.430 133.675 ;
        RECT 99.325 132.535 99.605 133.335 ;
        RECT 99.840 133.215 101.430 133.385 ;
        RECT 99.775 132.755 101.430 133.045 ;
        RECT 101.665 132.535 101.875 133.675 ;
        RECT 102.045 132.705 102.375 133.685 ;
        RECT 103.445 133.675 103.615 134.410 ;
        RECT 103.885 134.345 105.495 134.515 ;
        RECT 103.885 134.175 104.055 134.345 ;
        RECT 103.785 133.845 104.055 134.175 ;
        RECT 104.225 133.845 104.630 134.175 ;
        RECT 103.885 133.675 104.055 133.845 ;
        RECT 102.545 132.535 102.775 133.675 ;
        RECT 103.445 132.705 103.715 133.675 ;
        RECT 103.885 133.505 104.610 133.675 ;
        RECT 104.800 133.555 105.510 134.175 ;
        RECT 105.680 133.845 106.030 134.415 ;
        RECT 106.205 134.285 106.545 134.915 ;
        RECT 106.715 134.285 106.965 135.085 ;
        RECT 107.155 134.435 107.485 134.915 ;
        RECT 107.655 134.625 107.880 135.085 ;
        RECT 108.050 134.435 108.380 134.915 ;
        RECT 106.205 134.235 106.435 134.285 ;
        RECT 107.155 134.265 108.380 134.435 ;
        RECT 109.010 134.305 109.510 134.915 ;
        RECT 109.885 134.410 110.155 134.755 ;
        RECT 110.345 134.685 110.725 135.085 ;
        RECT 110.895 134.515 111.065 134.865 ;
        RECT 111.235 134.685 111.565 135.085 ;
        RECT 111.765 134.515 111.935 134.865 ;
        RECT 112.135 134.585 112.465 135.085 ;
        RECT 106.205 133.675 106.380 134.235 ;
        RECT 106.550 133.925 107.245 134.095 ;
        RECT 107.075 133.675 107.245 133.925 ;
        RECT 107.420 133.895 107.840 134.095 ;
        RECT 108.010 133.895 108.340 134.095 ;
        RECT 108.510 133.895 108.840 134.095 ;
        RECT 109.010 133.675 109.180 134.305 ;
        RECT 109.365 133.845 109.715 134.095 ;
        RECT 109.885 133.675 110.055 134.410 ;
        RECT 110.325 134.345 111.935 134.515 ;
        RECT 110.325 134.175 110.495 134.345 ;
        RECT 110.225 133.845 110.495 134.175 ;
        RECT 110.665 133.845 111.070 134.175 ;
        RECT 110.325 133.675 110.495 133.845 ;
        RECT 104.440 133.385 104.610 133.505 ;
        RECT 105.710 133.385 106.030 133.675 ;
        RECT 103.925 132.535 104.205 133.335 ;
        RECT 104.440 133.215 106.030 133.385 ;
        RECT 104.375 132.755 106.030 133.045 ;
        RECT 106.205 132.705 106.545 133.675 ;
        RECT 106.715 132.535 106.885 133.675 ;
        RECT 107.075 133.505 109.510 133.675 ;
        RECT 107.155 132.535 107.405 133.335 ;
        RECT 108.050 132.705 108.380 133.505 ;
        RECT 108.680 132.535 109.010 133.335 ;
        RECT 109.180 132.705 109.510 133.505 ;
        RECT 109.885 132.705 110.155 133.675 ;
        RECT 110.325 133.505 111.050 133.675 ;
        RECT 111.240 133.555 111.950 134.175 ;
        RECT 112.120 133.845 112.470 134.415 ;
        RECT 112.645 134.315 114.315 135.085 ;
        RECT 114.485 134.360 114.775 135.085 ;
        RECT 115.405 134.315 118.915 135.085 ;
        RECT 119.175 134.535 119.345 134.915 ;
        RECT 119.525 134.705 119.855 135.085 ;
        RECT 119.175 134.365 119.840 134.535 ;
        RECT 120.035 134.410 120.295 134.915 ;
        RECT 120.930 134.540 126.275 135.085 ;
        RECT 110.880 133.385 111.050 133.505 ;
        RECT 112.150 133.385 112.470 133.675 ;
        RECT 110.365 132.535 110.645 133.335 ;
        RECT 110.880 133.215 112.470 133.385 ;
        RECT 112.645 133.625 113.395 134.145 ;
        RECT 113.565 133.795 114.315 134.315 ;
        RECT 110.815 132.755 112.470 133.045 ;
        RECT 112.645 132.535 114.315 133.625 ;
        RECT 114.485 132.535 114.775 133.700 ;
        RECT 115.405 133.625 117.095 134.145 ;
        RECT 117.265 133.795 118.915 134.315 ;
        RECT 119.105 133.815 119.435 134.185 ;
        RECT 119.670 134.110 119.840 134.365 ;
        RECT 119.670 133.780 119.955 134.110 ;
        RECT 119.670 133.635 119.840 133.780 ;
        RECT 115.405 132.535 118.915 133.625 ;
        RECT 119.175 133.465 119.840 133.635 ;
        RECT 120.125 133.610 120.295 134.410 ;
        RECT 119.175 132.705 119.345 133.465 ;
        RECT 119.525 132.535 119.855 133.295 ;
        RECT 120.025 132.705 120.295 133.610 ;
        RECT 122.520 132.970 122.870 134.220 ;
        RECT 124.350 133.710 124.690 134.540 ;
        RECT 126.445 134.335 127.655 135.085 ;
        RECT 126.445 133.625 126.965 134.165 ;
        RECT 127.135 133.795 127.655 134.335 ;
        RECT 120.930 132.535 126.275 132.970 ;
        RECT 126.445 132.535 127.655 133.625 ;
        RECT 14.580 132.365 127.740 132.535 ;
        RECT 14.665 131.275 15.875 132.365 ;
        RECT 14.665 130.565 15.185 131.105 ;
        RECT 15.355 130.735 15.875 131.275 ;
        RECT 16.505 131.275 20.015 132.365 ;
        RECT 20.185 131.605 20.700 132.015 ;
        RECT 20.935 131.605 21.105 132.365 ;
        RECT 21.275 132.025 23.305 132.195 ;
        RECT 16.505 130.755 18.195 131.275 ;
        RECT 18.365 130.585 20.015 131.105 ;
        RECT 20.185 130.795 20.525 131.605 ;
        RECT 21.275 131.360 21.445 132.025 ;
        RECT 21.840 131.685 22.965 131.855 ;
        RECT 20.695 131.170 21.445 131.360 ;
        RECT 21.615 131.345 22.625 131.515 ;
        RECT 20.185 130.625 21.415 130.795 ;
        RECT 14.665 129.815 15.875 130.565 ;
        RECT 16.505 129.815 20.015 130.585 ;
        RECT 20.460 130.020 20.705 130.625 ;
        RECT 20.925 129.815 21.435 130.350 ;
        RECT 21.615 129.985 21.805 131.345 ;
        RECT 21.975 130.665 22.250 131.145 ;
        RECT 21.975 130.495 22.255 130.665 ;
        RECT 22.455 130.545 22.625 131.345 ;
        RECT 22.795 130.555 22.965 131.685 ;
        RECT 23.135 131.055 23.305 132.025 ;
        RECT 23.475 131.225 23.645 132.365 ;
        RECT 23.815 131.225 24.150 132.195 ;
        RECT 23.135 130.725 23.330 131.055 ;
        RECT 23.555 130.725 23.810 131.055 ;
        RECT 23.555 130.555 23.725 130.725 ;
        RECT 23.980 130.555 24.150 131.225 ;
        RECT 24.325 131.200 24.615 132.365 ;
        RECT 25.245 131.275 28.755 132.365 ;
        RECT 28.925 131.290 29.195 132.195 ;
        RECT 29.365 131.605 29.695 132.365 ;
        RECT 29.875 131.435 30.045 132.195 ;
        RECT 30.680 132.025 30.935 132.055 ;
        RECT 30.595 131.855 30.935 132.025 ;
        RECT 25.245 130.755 26.935 131.275 ;
        RECT 27.105 130.585 28.755 131.105 ;
        RECT 21.975 129.985 22.250 130.495 ;
        RECT 22.795 130.385 23.725 130.555 ;
        RECT 22.795 130.350 22.970 130.385 ;
        RECT 22.440 129.985 22.970 130.350 ;
        RECT 23.395 129.815 23.725 130.215 ;
        RECT 23.895 129.985 24.150 130.555 ;
        RECT 24.325 129.815 24.615 130.540 ;
        RECT 25.245 129.815 28.755 130.585 ;
        RECT 28.925 130.490 29.095 131.290 ;
        RECT 29.380 131.265 30.045 131.435 ;
        RECT 30.680 131.385 30.935 131.855 ;
        RECT 31.115 131.565 31.400 132.365 ;
        RECT 31.580 131.645 31.910 132.155 ;
        RECT 29.380 131.120 29.550 131.265 ;
        RECT 29.265 130.790 29.550 131.120 ;
        RECT 29.380 130.535 29.550 130.790 ;
        RECT 29.785 130.715 30.115 131.085 ;
        RECT 28.925 129.985 29.185 130.490 ;
        RECT 29.380 130.365 30.045 130.535 ;
        RECT 29.365 129.815 29.695 130.195 ;
        RECT 29.875 129.985 30.045 130.365 ;
        RECT 30.680 130.525 30.860 131.385 ;
        RECT 31.580 131.055 31.830 131.645 ;
        RECT 32.180 131.495 32.350 132.105 ;
        RECT 32.520 131.675 32.850 132.365 ;
        RECT 33.080 131.815 33.320 132.105 ;
        RECT 33.520 131.985 33.940 132.365 ;
        RECT 34.120 131.895 34.750 132.145 ;
        RECT 35.220 131.985 35.550 132.365 ;
        RECT 34.120 131.815 34.290 131.895 ;
        RECT 35.720 131.815 35.890 132.105 ;
        RECT 36.070 131.985 36.450 132.365 ;
        RECT 36.690 131.980 37.520 132.150 ;
        RECT 33.080 131.645 34.290 131.815 ;
        RECT 31.030 130.725 31.830 131.055 ;
        RECT 30.680 129.995 30.935 130.525 ;
        RECT 31.115 129.815 31.400 130.275 ;
        RECT 31.580 130.075 31.830 130.725 ;
        RECT 32.030 131.475 32.350 131.495 ;
        RECT 32.030 131.305 33.950 131.475 ;
        RECT 32.030 130.410 32.220 131.305 ;
        RECT 34.120 131.135 34.290 131.645 ;
        RECT 34.460 131.385 34.980 131.695 ;
        RECT 32.390 130.965 34.290 131.135 ;
        RECT 32.390 130.905 32.720 130.965 ;
        RECT 32.870 130.735 33.200 130.795 ;
        RECT 32.540 130.465 33.200 130.735 ;
        RECT 32.030 130.080 32.350 130.410 ;
        RECT 32.530 129.815 33.190 130.295 ;
        RECT 33.390 130.205 33.560 130.965 ;
        RECT 34.460 130.795 34.640 131.205 ;
        RECT 33.730 130.625 34.060 130.745 ;
        RECT 34.810 130.625 34.980 131.385 ;
        RECT 33.730 130.455 34.980 130.625 ;
        RECT 35.150 131.565 36.520 131.815 ;
        RECT 35.150 130.795 35.340 131.565 ;
        RECT 36.270 131.305 36.520 131.565 ;
        RECT 35.510 131.135 35.760 131.295 ;
        RECT 36.690 131.135 36.860 131.980 ;
        RECT 37.755 131.695 37.925 132.195 ;
        RECT 38.095 131.865 38.425 132.365 ;
        RECT 37.030 131.305 37.530 131.685 ;
        RECT 37.755 131.525 38.450 131.695 ;
        RECT 35.510 130.965 36.860 131.135 ;
        RECT 36.440 130.925 36.860 130.965 ;
        RECT 35.150 130.455 35.570 130.795 ;
        RECT 35.860 130.465 36.270 130.795 ;
        RECT 33.390 130.035 34.240 130.205 ;
        RECT 34.800 129.815 35.120 130.275 ;
        RECT 35.320 130.025 35.570 130.455 ;
        RECT 35.860 129.815 36.270 130.255 ;
        RECT 36.440 130.195 36.610 130.925 ;
        RECT 36.780 130.375 37.130 130.745 ;
        RECT 37.310 130.435 37.530 131.305 ;
        RECT 37.700 130.735 38.110 131.355 ;
        RECT 38.280 130.555 38.450 131.525 ;
        RECT 37.755 130.365 38.450 130.555 ;
        RECT 36.440 129.995 37.455 130.195 ;
        RECT 37.755 130.035 37.925 130.365 ;
        RECT 38.095 129.815 38.425 130.195 ;
        RECT 38.640 130.075 38.865 132.195 ;
        RECT 39.035 131.865 39.365 132.365 ;
        RECT 39.535 131.695 39.705 132.195 ;
        RECT 39.040 131.525 39.705 131.695 ;
        RECT 40.055 131.620 40.325 132.365 ;
        RECT 40.955 132.360 47.230 132.365 ;
        RECT 39.040 130.535 39.270 131.525 ;
        RECT 40.495 131.450 40.785 132.190 ;
        RECT 40.955 131.635 41.210 132.360 ;
        RECT 41.395 131.465 41.655 132.190 ;
        RECT 41.825 131.635 42.070 132.360 ;
        RECT 42.255 131.465 42.515 132.190 ;
        RECT 42.685 131.635 42.930 132.360 ;
        RECT 43.115 131.465 43.375 132.190 ;
        RECT 43.545 131.635 43.790 132.360 ;
        RECT 43.960 131.465 44.220 132.190 ;
        RECT 44.390 131.635 44.650 132.360 ;
        RECT 44.820 131.465 45.080 132.190 ;
        RECT 45.250 131.635 45.510 132.360 ;
        RECT 45.680 131.465 45.940 132.190 ;
        RECT 46.110 131.635 46.370 132.360 ;
        RECT 46.540 131.465 46.800 132.190 ;
        RECT 46.970 131.565 47.230 132.360 ;
        RECT 41.395 131.450 46.800 131.465 ;
        RECT 39.440 130.705 39.790 131.355 ;
        RECT 40.055 131.225 46.800 131.450 ;
        RECT 40.055 130.635 41.220 131.225 ;
        RECT 47.400 131.055 47.650 132.190 ;
        RECT 47.830 131.555 48.090 132.365 ;
        RECT 48.265 131.055 48.510 132.195 ;
        RECT 48.690 131.555 48.985 132.365 ;
        RECT 50.085 131.200 50.375 132.365 ;
        RECT 51.005 131.275 54.515 132.365 ;
        RECT 54.690 131.930 60.035 132.365 ;
        RECT 60.210 131.930 65.555 132.365 ;
        RECT 41.390 130.805 48.510 131.055 ;
        RECT 39.040 130.365 39.705 130.535 ;
        RECT 40.055 130.465 46.800 130.635 ;
        RECT 39.035 129.815 39.365 130.195 ;
        RECT 39.535 130.075 39.705 130.365 ;
        RECT 40.055 129.815 40.355 130.295 ;
        RECT 40.525 130.010 40.785 130.465 ;
        RECT 40.955 129.815 41.215 130.295 ;
        RECT 41.395 130.010 41.655 130.465 ;
        RECT 41.825 129.815 42.075 130.295 ;
        RECT 42.255 130.010 42.515 130.465 ;
        RECT 42.685 129.815 42.935 130.295 ;
        RECT 43.115 130.010 43.375 130.465 ;
        RECT 43.545 129.815 43.790 130.295 ;
        RECT 43.960 130.010 44.235 130.465 ;
        RECT 44.405 129.815 44.650 130.295 ;
        RECT 44.820 130.010 45.080 130.465 ;
        RECT 45.250 129.815 45.510 130.295 ;
        RECT 45.680 130.010 45.940 130.465 ;
        RECT 46.110 129.815 46.370 130.295 ;
        RECT 46.540 130.010 46.800 130.465 ;
        RECT 46.970 129.815 47.230 130.375 ;
        RECT 47.400 129.995 47.650 130.805 ;
        RECT 47.830 129.815 48.090 130.340 ;
        RECT 48.260 129.995 48.510 130.805 ;
        RECT 48.680 130.495 48.995 131.055 ;
        RECT 51.005 130.755 52.695 131.275 ;
        RECT 52.865 130.585 54.515 131.105 ;
        RECT 56.280 130.680 56.630 131.930 ;
        RECT 48.690 129.815 48.995 130.325 ;
        RECT 50.085 129.815 50.375 130.540 ;
        RECT 51.005 129.815 54.515 130.585 ;
        RECT 58.110 130.360 58.450 131.190 ;
        RECT 61.800 130.680 62.150 131.930 ;
        RECT 65.725 131.605 66.240 132.015 ;
        RECT 66.475 131.605 66.645 132.365 ;
        RECT 66.815 132.025 68.845 132.195 ;
        RECT 63.630 130.360 63.970 131.190 ;
        RECT 65.725 130.795 66.065 131.605 ;
        RECT 66.815 131.360 66.985 132.025 ;
        RECT 67.380 131.685 68.505 131.855 ;
        RECT 66.235 131.170 66.985 131.360 ;
        RECT 67.155 131.345 68.165 131.515 ;
        RECT 65.725 130.625 66.955 130.795 ;
        RECT 54.690 129.815 60.035 130.360 ;
        RECT 60.210 129.815 65.555 130.360 ;
        RECT 66.000 130.020 66.245 130.625 ;
        RECT 66.465 129.815 66.975 130.350 ;
        RECT 67.155 129.985 67.345 131.345 ;
        RECT 67.515 130.665 67.790 131.145 ;
        RECT 67.515 130.495 67.795 130.665 ;
        RECT 67.995 130.545 68.165 131.345 ;
        RECT 68.335 130.555 68.505 131.685 ;
        RECT 68.675 131.055 68.845 132.025 ;
        RECT 69.015 131.225 69.185 132.365 ;
        RECT 69.355 131.225 69.690 132.195 ;
        RECT 69.870 131.940 70.205 132.365 ;
        RECT 70.375 131.760 70.560 132.165 ;
        RECT 68.675 130.725 68.870 131.055 ;
        RECT 69.095 130.725 69.350 131.055 ;
        RECT 69.095 130.555 69.265 130.725 ;
        RECT 69.520 130.555 69.690 131.225 ;
        RECT 67.515 129.985 67.790 130.495 ;
        RECT 68.335 130.385 69.265 130.555 ;
        RECT 68.335 130.350 68.510 130.385 ;
        RECT 67.980 129.985 68.510 130.350 ;
        RECT 68.935 129.815 69.265 130.215 ;
        RECT 69.435 129.985 69.690 130.555 ;
        RECT 69.895 131.585 70.560 131.760 ;
        RECT 70.765 131.585 71.095 132.365 ;
        RECT 69.895 130.555 70.235 131.585 ;
        RECT 71.265 131.395 71.535 132.165 ;
        RECT 70.405 131.225 71.535 131.395 ;
        RECT 70.405 130.725 70.655 131.225 ;
        RECT 69.895 130.385 70.580 130.555 ;
        RECT 70.835 130.475 71.195 131.055 ;
        RECT 69.870 129.815 70.205 130.215 ;
        RECT 70.375 129.985 70.580 130.385 ;
        RECT 71.365 130.315 71.535 131.225 ;
        RECT 70.790 129.815 71.065 130.295 ;
        RECT 71.275 129.985 71.535 130.315 ;
        RECT 71.705 131.645 72.165 132.195 ;
        RECT 72.355 131.645 72.685 132.365 ;
        RECT 71.705 130.275 71.955 131.645 ;
        RECT 72.885 131.475 73.185 132.025 ;
        RECT 73.355 131.695 73.635 132.365 ;
        RECT 72.245 131.305 73.185 131.475 ;
        RECT 72.245 131.055 72.415 131.305 ;
        RECT 73.555 131.055 73.820 131.415 ;
        RECT 72.125 130.725 72.415 131.055 ;
        RECT 72.585 130.805 72.925 131.055 ;
        RECT 73.145 130.805 73.820 131.055 ;
        RECT 74.005 131.395 74.275 132.165 ;
        RECT 74.445 131.585 74.775 132.365 ;
        RECT 74.980 131.760 75.165 132.165 ;
        RECT 75.335 131.940 75.670 132.365 ;
        RECT 74.980 131.585 75.645 131.760 ;
        RECT 74.005 131.225 75.135 131.395 ;
        RECT 72.245 130.635 72.415 130.725 ;
        RECT 72.245 130.445 73.635 130.635 ;
        RECT 71.705 129.985 72.265 130.275 ;
        RECT 72.435 129.815 72.685 130.275 ;
        RECT 73.305 130.085 73.635 130.445 ;
        RECT 74.005 130.315 74.175 131.225 ;
        RECT 74.345 130.475 74.705 131.055 ;
        RECT 74.885 130.725 75.135 131.225 ;
        RECT 75.305 130.555 75.645 131.585 ;
        RECT 75.845 131.200 76.135 132.365 ;
        RECT 76.765 131.275 78.435 132.365 ;
        RECT 78.605 131.645 79.065 132.195 ;
        RECT 79.255 131.645 79.585 132.365 ;
        RECT 76.765 130.755 77.515 131.275 ;
        RECT 77.685 130.585 78.435 131.105 ;
        RECT 74.960 130.385 75.645 130.555 ;
        RECT 74.005 129.985 74.265 130.315 ;
        RECT 74.475 129.815 74.750 130.295 ;
        RECT 74.960 129.985 75.165 130.385 ;
        RECT 75.335 129.815 75.670 130.215 ;
        RECT 75.845 129.815 76.135 130.540 ;
        RECT 76.765 129.815 78.435 130.585 ;
        RECT 78.605 130.275 78.855 131.645 ;
        RECT 79.785 131.475 80.085 132.025 ;
        RECT 80.255 131.695 80.535 132.365 ;
        RECT 79.145 131.305 80.085 131.475 ;
        RECT 79.145 131.055 79.315 131.305 ;
        RECT 80.455 131.055 80.720 131.415 ;
        RECT 79.025 130.725 79.315 131.055 ;
        RECT 79.485 130.805 79.825 131.055 ;
        RECT 80.045 130.805 80.720 131.055 ;
        RECT 80.905 131.275 83.495 132.365 ;
        RECT 83.670 131.930 89.015 132.365 ;
        RECT 80.905 130.755 82.115 131.275 ;
        RECT 79.145 130.635 79.315 130.725 ;
        RECT 79.145 130.445 80.535 130.635 ;
        RECT 82.285 130.585 83.495 131.105 ;
        RECT 85.260 130.680 85.610 131.930 ;
        RECT 89.225 131.225 89.455 132.365 ;
        RECT 89.625 131.215 89.955 132.195 ;
        RECT 90.125 131.225 90.335 132.365 ;
        RECT 90.675 131.565 90.845 132.365 ;
        RECT 91.015 131.345 91.345 132.195 ;
        RECT 91.515 131.565 91.685 132.365 ;
        RECT 91.855 131.345 92.185 132.195 ;
        RECT 92.355 131.565 92.525 132.365 ;
        RECT 92.695 131.345 93.025 132.195 ;
        RECT 93.195 131.565 93.365 132.365 ;
        RECT 93.535 131.345 93.865 132.195 ;
        RECT 94.035 131.565 94.205 132.365 ;
        RECT 94.375 131.345 94.705 132.195 ;
        RECT 94.875 131.565 95.045 132.365 ;
        RECT 95.215 131.345 95.545 132.195 ;
        RECT 95.715 131.565 95.885 132.365 ;
        RECT 96.055 131.345 96.385 132.195 ;
        RECT 96.555 131.565 96.725 132.365 ;
        RECT 96.895 131.345 97.225 132.195 ;
        RECT 97.395 131.565 97.565 132.365 ;
        RECT 97.735 131.345 98.065 132.195 ;
        RECT 98.235 131.565 98.405 132.365 ;
        RECT 98.575 131.345 98.905 132.195 ;
        RECT 99.075 131.565 99.245 132.365 ;
        RECT 99.415 131.345 99.745 132.195 ;
        RECT 99.915 131.515 100.085 132.365 ;
        RECT 100.255 131.345 100.585 132.195 ;
        RECT 100.755 131.515 100.925 132.365 ;
        RECT 101.095 131.345 101.425 132.195 ;
        RECT 78.605 129.985 79.165 130.275 ;
        RECT 79.335 129.815 79.585 130.275 ;
        RECT 80.205 130.085 80.535 130.445 ;
        RECT 80.905 129.815 83.495 130.585 ;
        RECT 87.090 130.360 87.430 131.190 ;
        RECT 89.205 130.805 89.535 131.055 ;
        RECT 83.670 129.815 89.015 130.360 ;
        RECT 89.225 129.815 89.455 130.635 ;
        RECT 89.705 130.615 89.955 131.215 ;
        RECT 90.565 131.175 97.225 131.345 ;
        RECT 97.395 131.175 99.745 131.345 ;
        RECT 99.915 131.175 101.425 131.345 ;
        RECT 101.605 131.200 101.895 132.365 ;
        RECT 102.525 131.275 104.195 132.365 ;
        RECT 104.370 131.930 109.715 132.365 ;
        RECT 90.565 130.635 90.840 131.175 ;
        RECT 97.395 131.005 97.570 131.175 ;
        RECT 99.915 131.005 100.085 131.175 ;
        RECT 91.010 130.805 97.570 131.005 ;
        RECT 97.775 130.805 100.085 131.005 ;
        RECT 100.255 130.805 101.430 131.005 ;
        RECT 97.395 130.635 97.570 130.805 ;
        RECT 99.915 130.635 100.085 130.805 ;
        RECT 102.525 130.755 103.275 131.275 ;
        RECT 89.625 129.985 89.955 130.615 ;
        RECT 90.125 129.815 90.335 130.635 ;
        RECT 90.565 130.465 97.225 130.635 ;
        RECT 97.395 130.465 99.745 130.635 ;
        RECT 99.915 130.465 101.425 130.635 ;
        RECT 103.445 130.585 104.195 131.105 ;
        RECT 105.960 130.680 106.310 131.930 ;
        RECT 109.885 131.645 110.345 132.195 ;
        RECT 110.535 131.645 110.865 132.365 ;
        RECT 90.675 129.815 90.845 130.295 ;
        RECT 91.015 129.990 91.345 130.465 ;
        RECT 91.515 129.815 91.685 130.295 ;
        RECT 91.855 129.990 92.185 130.465 ;
        RECT 92.355 129.815 92.525 130.295 ;
        RECT 92.695 129.990 93.025 130.465 ;
        RECT 93.195 129.815 93.365 130.295 ;
        RECT 93.535 129.990 93.865 130.465 ;
        RECT 94.035 129.815 94.205 130.295 ;
        RECT 94.375 129.990 94.705 130.465 ;
        RECT 94.875 129.815 95.045 130.295 ;
        RECT 95.215 129.990 95.545 130.465 ;
        RECT 95.295 129.985 95.465 129.990 ;
        RECT 95.715 129.815 95.885 130.295 ;
        RECT 96.055 129.990 96.385 130.465 ;
        RECT 96.135 129.985 96.305 129.990 ;
        RECT 96.555 129.815 96.725 130.295 ;
        RECT 96.895 129.990 97.225 130.465 ;
        RECT 96.975 129.985 97.225 129.990 ;
        RECT 97.395 129.815 97.565 130.295 ;
        RECT 97.735 129.990 98.065 130.465 ;
        RECT 98.235 129.815 98.405 130.295 ;
        RECT 98.575 129.990 98.905 130.465 ;
        RECT 99.075 129.815 99.245 130.295 ;
        RECT 99.415 129.990 99.745 130.465 ;
        RECT 99.915 129.815 100.085 130.295 ;
        RECT 100.255 129.990 100.585 130.465 ;
        RECT 100.755 129.815 100.925 130.295 ;
        RECT 101.095 129.990 101.425 130.465 ;
        RECT 101.605 129.815 101.895 130.540 ;
        RECT 102.525 129.815 104.195 130.585 ;
        RECT 107.790 130.360 108.130 131.190 ;
        RECT 104.370 129.815 109.715 130.360 ;
        RECT 109.885 130.275 110.135 131.645 ;
        RECT 111.065 131.475 111.365 132.025 ;
        RECT 111.535 131.695 111.815 132.365 ;
        RECT 110.425 131.305 111.365 131.475 ;
        RECT 110.425 131.055 110.595 131.305 ;
        RECT 111.735 131.055 112.000 131.415 ;
        RECT 110.305 130.725 110.595 131.055 ;
        RECT 110.765 130.805 111.105 131.055 ;
        RECT 111.325 130.805 112.000 131.055 ;
        RECT 112.645 131.275 115.235 132.365 ;
        RECT 115.410 131.930 120.755 132.365 ;
        RECT 120.930 131.930 126.275 132.365 ;
        RECT 112.645 130.755 113.855 131.275 ;
        RECT 110.425 130.635 110.595 130.725 ;
        RECT 110.425 130.445 111.815 130.635 ;
        RECT 114.025 130.585 115.235 131.105 ;
        RECT 117.000 130.680 117.350 131.930 ;
        RECT 109.885 129.985 110.445 130.275 ;
        RECT 110.615 129.815 110.865 130.275 ;
        RECT 111.485 130.085 111.815 130.445 ;
        RECT 112.645 129.815 115.235 130.585 ;
        RECT 118.830 130.360 119.170 131.190 ;
        RECT 122.520 130.680 122.870 131.930 ;
        RECT 126.445 131.275 127.655 132.365 ;
        RECT 124.350 130.360 124.690 131.190 ;
        RECT 126.445 130.735 126.965 131.275 ;
        RECT 127.135 130.565 127.655 131.105 ;
        RECT 115.410 129.815 120.755 130.360 ;
        RECT 120.930 129.815 126.275 130.360 ;
        RECT 126.445 129.815 127.655 130.565 ;
        RECT 14.580 129.645 127.740 129.815 ;
        RECT 14.665 128.895 15.875 129.645 ;
        RECT 16.045 128.895 17.255 129.645 ;
        RECT 17.800 129.305 18.055 129.465 ;
        RECT 17.715 129.135 18.055 129.305 ;
        RECT 18.235 129.185 18.520 129.645 ;
        RECT 14.665 128.355 15.185 128.895 ;
        RECT 15.355 128.185 15.875 128.725 ;
        RECT 14.665 127.095 15.875 128.185 ;
        RECT 16.045 128.185 16.565 128.725 ;
        RECT 16.735 128.355 17.255 128.895 ;
        RECT 17.800 128.935 18.055 129.135 ;
        RECT 16.045 127.095 17.255 128.185 ;
        RECT 17.800 128.075 17.980 128.935 ;
        RECT 18.700 128.735 18.950 129.385 ;
        RECT 18.150 128.405 18.950 128.735 ;
        RECT 17.800 127.405 18.055 128.075 ;
        RECT 18.235 127.095 18.520 127.895 ;
        RECT 18.700 127.815 18.950 128.405 ;
        RECT 19.150 129.050 19.470 129.380 ;
        RECT 19.650 129.165 20.310 129.645 ;
        RECT 20.510 129.255 21.360 129.425 ;
        RECT 19.150 128.155 19.340 129.050 ;
        RECT 19.660 128.725 20.320 128.995 ;
        RECT 19.990 128.665 20.320 128.725 ;
        RECT 19.510 128.495 19.840 128.555 ;
        RECT 20.510 128.495 20.680 129.255 ;
        RECT 21.920 129.185 22.240 129.645 ;
        RECT 22.440 129.005 22.690 129.435 ;
        RECT 22.980 129.205 23.390 129.645 ;
        RECT 23.560 129.265 24.575 129.465 ;
        RECT 20.850 128.835 22.100 129.005 ;
        RECT 20.850 128.715 21.180 128.835 ;
        RECT 19.510 128.325 21.410 128.495 ;
        RECT 19.150 127.985 21.070 128.155 ;
        RECT 19.150 127.965 19.470 127.985 ;
        RECT 18.700 127.305 19.030 127.815 ;
        RECT 19.300 127.355 19.470 127.965 ;
        RECT 21.240 127.815 21.410 128.325 ;
        RECT 21.580 128.255 21.760 128.665 ;
        RECT 21.930 128.075 22.100 128.835 ;
        RECT 19.640 127.095 19.970 127.785 ;
        RECT 20.200 127.645 21.410 127.815 ;
        RECT 21.580 127.765 22.100 128.075 ;
        RECT 22.270 128.665 22.690 129.005 ;
        RECT 22.980 128.665 23.390 128.995 ;
        RECT 22.270 127.895 22.460 128.665 ;
        RECT 23.560 128.535 23.730 129.265 ;
        RECT 24.875 129.095 25.045 129.425 ;
        RECT 25.215 129.265 25.545 129.645 ;
        RECT 23.900 128.715 24.250 129.085 ;
        RECT 23.560 128.495 23.980 128.535 ;
        RECT 22.630 128.325 23.980 128.495 ;
        RECT 22.630 128.165 22.880 128.325 ;
        RECT 23.390 127.895 23.640 128.155 ;
        RECT 22.270 127.645 23.640 127.895 ;
        RECT 20.200 127.355 20.440 127.645 ;
        RECT 21.240 127.565 21.410 127.645 ;
        RECT 20.640 127.095 21.060 127.475 ;
        RECT 21.240 127.315 21.870 127.565 ;
        RECT 22.340 127.095 22.670 127.475 ;
        RECT 22.840 127.355 23.010 127.645 ;
        RECT 23.810 127.480 23.980 128.325 ;
        RECT 24.430 128.155 24.650 129.025 ;
        RECT 24.875 128.905 25.570 129.095 ;
        RECT 24.150 127.775 24.650 128.155 ;
        RECT 24.820 128.105 25.230 128.725 ;
        RECT 25.400 127.935 25.570 128.905 ;
        RECT 24.875 127.765 25.570 127.935 ;
        RECT 23.190 127.095 23.570 127.475 ;
        RECT 23.810 127.310 24.640 127.480 ;
        RECT 24.875 127.265 25.045 127.765 ;
        RECT 25.215 127.095 25.545 127.595 ;
        RECT 25.760 127.265 25.985 129.385 ;
        RECT 26.155 129.265 26.485 129.645 ;
        RECT 26.655 129.095 26.825 129.385 ;
        RECT 28.010 129.100 33.355 129.645 ;
        RECT 26.160 128.925 26.825 129.095 ;
        RECT 26.160 127.935 26.390 128.925 ;
        RECT 26.560 128.105 26.910 128.755 ;
        RECT 26.160 127.765 26.825 127.935 ;
        RECT 26.155 127.095 26.485 127.595 ;
        RECT 26.655 127.265 26.825 127.765 ;
        RECT 29.600 127.530 29.950 128.780 ;
        RECT 31.430 128.270 31.770 129.100 ;
        RECT 33.565 128.825 33.795 129.645 ;
        RECT 33.965 128.845 34.295 129.475 ;
        RECT 33.545 128.405 33.875 128.655 ;
        RECT 34.045 128.245 34.295 128.845 ;
        RECT 34.465 128.825 34.675 129.645 ;
        RECT 35.365 128.875 37.035 129.645 ;
        RECT 37.205 128.920 37.495 129.645 ;
        RECT 38.585 128.970 38.845 129.475 ;
        RECT 39.025 129.265 39.355 129.645 ;
        RECT 39.535 129.095 39.705 129.475 ;
        RECT 28.010 127.095 33.355 127.530 ;
        RECT 33.565 127.095 33.795 128.235 ;
        RECT 33.965 127.265 34.295 128.245 ;
        RECT 34.465 127.095 34.675 128.235 ;
        RECT 35.365 128.185 36.115 128.705 ;
        RECT 36.285 128.355 37.035 128.875 ;
        RECT 35.365 127.095 37.035 128.185 ;
        RECT 37.205 127.095 37.495 128.260 ;
        RECT 38.585 128.170 38.755 128.970 ;
        RECT 39.040 128.925 39.705 129.095 ;
        RECT 40.165 129.015 40.495 129.375 ;
        RECT 41.115 129.185 41.365 129.645 ;
        RECT 41.535 129.185 42.095 129.475 ;
        RECT 39.040 128.670 39.210 128.925 ;
        RECT 40.165 128.825 41.555 129.015 ;
        RECT 38.925 128.340 39.210 128.670 ;
        RECT 39.445 128.375 39.775 128.745 ;
        RECT 41.385 128.735 41.555 128.825 ;
        RECT 39.980 128.405 40.655 128.655 ;
        RECT 40.875 128.405 41.215 128.655 ;
        RECT 41.385 128.405 41.675 128.735 ;
        RECT 39.040 128.195 39.210 128.340 ;
        RECT 38.585 127.265 38.855 128.170 ;
        RECT 39.040 128.025 39.705 128.195 ;
        RECT 39.980 128.045 40.245 128.405 ;
        RECT 41.385 128.155 41.555 128.405 ;
        RECT 39.025 127.095 39.355 127.855 ;
        RECT 39.535 127.265 39.705 128.025 ;
        RECT 40.615 127.985 41.555 128.155 ;
        RECT 40.165 127.095 40.445 127.765 ;
        RECT 40.615 127.435 40.915 127.985 ;
        RECT 41.845 127.815 42.095 129.185 ;
        RECT 42.465 129.015 42.795 129.375 ;
        RECT 43.415 129.185 43.665 129.645 ;
        RECT 43.835 129.185 44.395 129.475 ;
        RECT 42.465 128.825 43.855 129.015 ;
        RECT 43.685 128.735 43.855 128.825 ;
        RECT 42.280 128.405 42.955 128.655 ;
        RECT 43.175 128.405 43.515 128.655 ;
        RECT 43.685 128.405 43.975 128.735 ;
        RECT 42.280 128.045 42.545 128.405 ;
        RECT 43.685 128.155 43.855 128.405 ;
        RECT 41.115 127.095 41.445 127.815 ;
        RECT 41.635 127.265 42.095 127.815 ;
        RECT 42.915 127.985 43.855 128.155 ;
        RECT 42.465 127.095 42.745 127.765 ;
        RECT 42.915 127.435 43.215 127.985 ;
        RECT 44.145 127.815 44.395 129.185 ;
        RECT 45.235 128.955 45.565 129.645 ;
        RECT 46.025 129.050 46.645 129.475 ;
        RECT 46.815 129.155 47.145 129.645 ;
        RECT 46.285 128.715 46.645 129.050 ;
        RECT 47.525 129.015 47.855 129.375 ;
        RECT 48.475 129.185 48.725 129.645 ;
        RECT 48.895 129.185 49.455 129.475 ;
        RECT 45.225 128.435 46.645 128.715 ;
        RECT 43.415 127.095 43.745 127.815 ;
        RECT 43.935 127.265 44.395 127.815 ;
        RECT 44.695 127.095 45.025 128.265 ;
        RECT 45.225 127.265 45.555 128.435 ;
        RECT 45.755 127.095 46.085 128.265 ;
        RECT 46.285 127.265 46.645 128.435 ;
        RECT 46.815 128.405 47.155 128.985 ;
        RECT 47.525 128.825 48.915 129.015 ;
        RECT 48.745 128.735 48.915 128.825 ;
        RECT 47.340 128.405 48.015 128.655 ;
        RECT 48.235 128.405 48.575 128.655 ;
        RECT 48.745 128.405 49.035 128.735 ;
        RECT 46.815 127.095 47.145 128.235 ;
        RECT 47.340 128.045 47.605 128.405 ;
        RECT 48.745 128.155 48.915 128.405 ;
        RECT 47.975 127.985 48.915 128.155 ;
        RECT 47.525 127.095 47.805 127.765 ;
        RECT 47.975 127.435 48.275 127.985 ;
        RECT 49.205 127.815 49.455 129.185 ;
        RECT 49.625 128.895 50.835 129.645 ;
        RECT 48.475 127.095 48.805 127.815 ;
        RECT 48.995 127.265 49.455 127.815 ;
        RECT 49.625 128.185 50.145 128.725 ;
        RECT 50.315 128.355 50.835 128.895 ;
        RECT 51.005 128.875 54.515 129.645 ;
        RECT 51.005 128.185 52.695 128.705 ;
        RECT 52.865 128.355 54.515 128.875 ;
        RECT 54.960 128.835 55.205 129.440 ;
        RECT 55.425 129.110 55.935 129.645 ;
        RECT 54.685 128.665 55.915 128.835 ;
        RECT 49.625 127.095 50.835 128.185 ;
        RECT 51.005 127.095 54.515 128.185 ;
        RECT 54.685 127.855 55.025 128.665 ;
        RECT 55.195 128.100 55.945 128.290 ;
        RECT 54.685 127.445 55.200 127.855 ;
        RECT 55.435 127.095 55.605 127.855 ;
        RECT 55.775 127.435 55.945 128.100 ;
        RECT 56.115 128.115 56.305 129.475 ;
        RECT 56.475 129.305 56.750 129.475 ;
        RECT 56.475 129.135 56.755 129.305 ;
        RECT 56.475 128.315 56.750 129.135 ;
        RECT 56.940 129.110 57.470 129.475 ;
        RECT 57.895 129.245 58.225 129.645 ;
        RECT 57.295 129.075 57.470 129.110 ;
        RECT 56.955 128.115 57.125 128.915 ;
        RECT 56.115 127.945 57.125 128.115 ;
        RECT 57.295 128.905 58.225 129.075 ;
        RECT 58.395 128.905 58.650 129.475 ;
        RECT 57.295 127.775 57.465 128.905 ;
        RECT 58.055 128.735 58.225 128.905 ;
        RECT 56.340 127.605 57.465 127.775 ;
        RECT 57.635 128.405 57.830 128.735 ;
        RECT 58.055 128.405 58.310 128.735 ;
        RECT 57.635 127.435 57.805 128.405 ;
        RECT 58.480 128.235 58.650 128.905 ;
        RECT 59.285 128.875 62.795 129.645 ;
        RECT 62.965 128.920 63.255 129.645 ;
        RECT 63.425 128.895 64.635 129.645 ;
        RECT 65.180 129.305 65.435 129.465 ;
        RECT 65.095 129.135 65.435 129.305 ;
        RECT 65.615 129.185 65.900 129.645 ;
        RECT 55.775 127.265 57.805 127.435 ;
        RECT 57.975 127.095 58.145 128.235 ;
        RECT 58.315 127.265 58.650 128.235 ;
        RECT 59.285 128.185 60.975 128.705 ;
        RECT 61.145 128.355 62.795 128.875 ;
        RECT 59.285 127.095 62.795 128.185 ;
        RECT 62.965 127.095 63.255 128.260 ;
        RECT 63.425 128.185 63.945 128.725 ;
        RECT 64.115 128.355 64.635 128.895 ;
        RECT 65.180 128.935 65.435 129.135 ;
        RECT 63.425 127.095 64.635 128.185 ;
        RECT 65.180 128.075 65.360 128.935 ;
        RECT 66.080 128.735 66.330 129.385 ;
        RECT 65.530 128.405 66.330 128.735 ;
        RECT 65.180 127.405 65.435 128.075 ;
        RECT 65.615 127.095 65.900 127.895 ;
        RECT 66.080 127.815 66.330 128.405 ;
        RECT 66.530 129.050 66.850 129.380 ;
        RECT 67.030 129.165 67.690 129.645 ;
        RECT 67.890 129.255 68.740 129.425 ;
        RECT 66.530 128.155 66.720 129.050 ;
        RECT 67.040 128.725 67.700 128.995 ;
        RECT 67.370 128.665 67.700 128.725 ;
        RECT 66.890 128.495 67.220 128.555 ;
        RECT 67.890 128.495 68.060 129.255 ;
        RECT 69.300 129.185 69.620 129.645 ;
        RECT 69.820 129.005 70.070 129.435 ;
        RECT 70.360 129.205 70.770 129.645 ;
        RECT 70.940 129.265 71.955 129.465 ;
        RECT 68.230 128.835 69.480 129.005 ;
        RECT 68.230 128.715 68.560 128.835 ;
        RECT 66.890 128.325 68.790 128.495 ;
        RECT 66.530 127.985 68.450 128.155 ;
        RECT 66.530 127.965 66.850 127.985 ;
        RECT 66.080 127.305 66.410 127.815 ;
        RECT 66.680 127.355 66.850 127.965 ;
        RECT 68.620 127.815 68.790 128.325 ;
        RECT 68.960 128.255 69.140 128.665 ;
        RECT 69.310 128.075 69.480 128.835 ;
        RECT 67.020 127.095 67.350 127.785 ;
        RECT 67.580 127.645 68.790 127.815 ;
        RECT 68.960 127.765 69.480 128.075 ;
        RECT 69.650 128.665 70.070 129.005 ;
        RECT 70.360 128.665 70.770 128.995 ;
        RECT 69.650 127.895 69.840 128.665 ;
        RECT 70.940 128.535 71.110 129.265 ;
        RECT 72.255 129.095 72.425 129.425 ;
        RECT 72.595 129.265 72.925 129.645 ;
        RECT 71.280 128.715 71.630 129.085 ;
        RECT 70.940 128.495 71.360 128.535 ;
        RECT 70.010 128.325 71.360 128.495 ;
        RECT 70.010 128.165 70.260 128.325 ;
        RECT 70.770 127.895 71.020 128.155 ;
        RECT 69.650 127.645 71.020 127.895 ;
        RECT 67.580 127.355 67.820 127.645 ;
        RECT 68.620 127.565 68.790 127.645 ;
        RECT 68.020 127.095 68.440 127.475 ;
        RECT 68.620 127.315 69.250 127.565 ;
        RECT 69.720 127.095 70.050 127.475 ;
        RECT 70.220 127.355 70.390 127.645 ;
        RECT 71.190 127.480 71.360 128.325 ;
        RECT 71.810 128.155 72.030 129.025 ;
        RECT 72.255 128.905 72.950 129.095 ;
        RECT 71.530 127.775 72.030 128.155 ;
        RECT 72.200 128.105 72.610 128.725 ;
        RECT 72.780 127.935 72.950 128.905 ;
        RECT 72.255 127.765 72.950 127.935 ;
        RECT 70.570 127.095 70.950 127.475 ;
        RECT 71.190 127.310 72.020 127.480 ;
        RECT 72.255 127.265 72.425 127.765 ;
        RECT 72.595 127.095 72.925 127.595 ;
        RECT 73.140 127.265 73.365 129.385 ;
        RECT 73.535 129.265 73.865 129.645 ;
        RECT 74.035 129.095 74.205 129.385 ;
        RECT 73.540 128.925 74.205 129.095 ;
        RECT 74.665 129.015 74.995 129.375 ;
        RECT 75.615 129.185 75.865 129.645 ;
        RECT 76.035 129.185 76.595 129.475 ;
        RECT 73.540 127.935 73.770 128.925 ;
        RECT 74.665 128.825 76.055 129.015 ;
        RECT 73.940 128.105 74.290 128.755 ;
        RECT 75.885 128.735 76.055 128.825 ;
        RECT 74.480 128.405 75.155 128.655 ;
        RECT 75.375 128.405 75.715 128.655 ;
        RECT 75.885 128.405 76.175 128.735 ;
        RECT 74.480 128.045 74.745 128.405 ;
        RECT 75.885 128.155 76.055 128.405 ;
        RECT 75.115 127.985 76.055 128.155 ;
        RECT 73.540 127.765 74.205 127.935 ;
        RECT 73.535 127.095 73.865 127.595 ;
        RECT 74.035 127.265 74.205 127.765 ;
        RECT 74.665 127.095 74.945 127.765 ;
        RECT 75.115 127.435 75.415 127.985 ;
        RECT 76.345 127.815 76.595 129.185 ;
        RECT 76.965 129.015 77.295 129.375 ;
        RECT 77.915 129.185 78.165 129.645 ;
        RECT 78.335 129.185 78.895 129.475 ;
        RECT 76.965 128.825 78.355 129.015 ;
        RECT 78.185 128.735 78.355 128.825 ;
        RECT 76.780 128.405 77.455 128.655 ;
        RECT 77.675 128.405 78.015 128.655 ;
        RECT 78.185 128.405 78.475 128.735 ;
        RECT 76.780 128.045 77.045 128.405 ;
        RECT 78.185 128.155 78.355 128.405 ;
        RECT 75.615 127.095 75.945 127.815 ;
        RECT 76.135 127.265 76.595 127.815 ;
        RECT 77.415 127.985 78.355 128.155 ;
        RECT 76.965 127.095 77.245 127.765 ;
        RECT 77.415 127.435 77.715 127.985 ;
        RECT 78.645 127.815 78.895 129.185 ;
        RECT 79.340 128.835 79.585 129.440 ;
        RECT 79.805 129.110 80.315 129.645 ;
        RECT 77.915 127.095 78.245 127.815 ;
        RECT 78.435 127.265 78.895 127.815 ;
        RECT 79.065 128.665 80.295 128.835 ;
        RECT 79.065 127.855 79.405 128.665 ;
        RECT 79.575 128.100 80.325 128.290 ;
        RECT 79.065 127.445 79.580 127.855 ;
        RECT 79.815 127.095 79.985 127.855 ;
        RECT 80.155 127.435 80.325 128.100 ;
        RECT 80.495 128.115 80.685 129.475 ;
        RECT 80.855 128.625 81.130 129.475 ;
        RECT 81.320 129.110 81.850 129.475 ;
        RECT 82.275 129.245 82.605 129.645 ;
        RECT 81.675 129.075 81.850 129.110 ;
        RECT 80.855 128.455 81.135 128.625 ;
        RECT 80.855 128.315 81.130 128.455 ;
        RECT 81.335 128.115 81.505 128.915 ;
        RECT 80.495 127.945 81.505 128.115 ;
        RECT 81.675 128.905 82.605 129.075 ;
        RECT 82.775 128.905 83.030 129.475 ;
        RECT 81.675 127.775 81.845 128.905 ;
        RECT 82.435 128.735 82.605 128.905 ;
        RECT 80.720 127.605 81.845 127.775 ;
        RECT 82.015 128.405 82.210 128.735 ;
        RECT 82.435 128.405 82.690 128.735 ;
        RECT 82.015 127.435 82.185 128.405 ;
        RECT 82.860 128.235 83.030 128.905 ;
        RECT 80.155 127.265 82.185 127.435 ;
        RECT 82.355 127.095 82.525 128.235 ;
        RECT 82.695 127.265 83.030 128.235 ;
        RECT 83.205 129.185 83.765 129.475 ;
        RECT 83.935 129.185 84.185 129.645 ;
        RECT 83.205 127.815 83.455 129.185 ;
        RECT 84.805 129.015 85.135 129.375 ;
        RECT 83.745 128.825 85.135 129.015 ;
        RECT 85.505 128.875 87.175 129.645 ;
        RECT 87.435 129.095 87.605 129.475 ;
        RECT 87.785 129.265 88.115 129.645 ;
        RECT 87.435 128.925 88.100 129.095 ;
        RECT 88.295 128.970 88.555 129.475 ;
        RECT 83.745 128.735 83.915 128.825 ;
        RECT 83.625 128.405 83.915 128.735 ;
        RECT 84.085 128.405 84.425 128.655 ;
        RECT 84.645 128.405 85.320 128.655 ;
        RECT 83.745 128.155 83.915 128.405 ;
        RECT 83.745 127.985 84.685 128.155 ;
        RECT 85.055 128.045 85.320 128.405 ;
        RECT 85.505 128.185 86.255 128.705 ;
        RECT 86.425 128.355 87.175 128.875 ;
        RECT 87.365 128.375 87.695 128.745 ;
        RECT 87.930 128.670 88.100 128.925 ;
        RECT 87.930 128.340 88.215 128.670 ;
        RECT 87.930 128.195 88.100 128.340 ;
        RECT 83.205 127.265 83.665 127.815 ;
        RECT 83.855 127.095 84.185 127.815 ;
        RECT 84.385 127.435 84.685 127.985 ;
        RECT 84.855 127.095 85.135 127.765 ;
        RECT 85.505 127.095 87.175 128.185 ;
        RECT 87.435 128.025 88.100 128.195 ;
        RECT 88.385 128.170 88.555 128.970 ;
        RECT 88.725 128.920 89.015 129.645 ;
        RECT 89.650 128.905 89.905 129.475 ;
        RECT 90.075 129.245 90.405 129.645 ;
        RECT 90.830 129.110 91.360 129.475 ;
        RECT 90.830 129.075 91.005 129.110 ;
        RECT 90.075 128.905 91.005 129.075 ;
        RECT 87.435 127.265 87.605 128.025 ;
        RECT 87.785 127.095 88.115 127.855 ;
        RECT 88.285 127.265 88.555 128.170 ;
        RECT 88.725 127.095 89.015 128.260 ;
        RECT 89.650 128.235 89.820 128.905 ;
        RECT 90.075 128.735 90.245 128.905 ;
        RECT 89.990 128.405 90.245 128.735 ;
        RECT 90.470 128.405 90.665 128.735 ;
        RECT 89.650 127.265 89.985 128.235 ;
        RECT 90.155 127.095 90.325 128.235 ;
        RECT 90.495 127.435 90.665 128.405 ;
        RECT 90.835 127.775 91.005 128.905 ;
        RECT 91.175 128.115 91.345 128.915 ;
        RECT 91.550 128.625 91.825 129.475 ;
        RECT 91.545 128.455 91.825 128.625 ;
        RECT 91.550 128.315 91.825 128.455 ;
        RECT 91.995 128.115 92.185 129.475 ;
        RECT 92.365 129.110 92.875 129.645 ;
        RECT 93.095 128.835 93.340 129.440 ;
        RECT 94.335 129.095 94.505 129.475 ;
        RECT 94.685 129.265 95.015 129.645 ;
        RECT 94.335 128.925 95.000 129.095 ;
        RECT 95.195 128.970 95.455 129.475 ;
        RECT 95.625 129.135 95.930 129.645 ;
        RECT 92.385 128.665 93.615 128.835 ;
        RECT 91.175 127.945 92.185 128.115 ;
        RECT 92.355 128.100 93.105 128.290 ;
        RECT 90.835 127.605 91.960 127.775 ;
        RECT 92.355 127.435 92.525 128.100 ;
        RECT 93.275 127.855 93.615 128.665 ;
        RECT 94.265 128.375 94.595 128.745 ;
        RECT 94.830 128.670 95.000 128.925 ;
        RECT 94.830 128.340 95.115 128.670 ;
        RECT 94.830 128.195 95.000 128.340 ;
        RECT 90.495 127.265 92.525 127.435 ;
        RECT 92.695 127.095 92.865 127.855 ;
        RECT 93.100 127.445 93.615 127.855 ;
        RECT 94.335 128.025 95.000 128.195 ;
        RECT 95.285 128.170 95.455 128.970 ;
        RECT 95.625 128.405 95.940 128.965 ;
        RECT 96.110 128.655 96.360 129.465 ;
        RECT 96.530 129.120 96.790 129.645 ;
        RECT 96.970 128.655 97.220 129.465 ;
        RECT 97.390 129.085 97.650 129.645 ;
        RECT 97.820 128.995 98.080 129.450 ;
        RECT 98.250 129.165 98.510 129.645 ;
        RECT 98.680 128.995 98.940 129.450 ;
        RECT 99.110 129.165 99.370 129.645 ;
        RECT 99.540 128.995 99.800 129.450 ;
        RECT 99.970 129.165 100.215 129.645 ;
        RECT 100.385 128.995 100.660 129.450 ;
        RECT 100.830 129.165 101.075 129.645 ;
        RECT 101.245 128.995 101.505 129.450 ;
        RECT 101.685 129.165 101.935 129.645 ;
        RECT 102.105 128.995 102.365 129.450 ;
        RECT 102.545 129.165 102.795 129.645 ;
        RECT 102.965 128.995 103.225 129.450 ;
        RECT 103.405 129.165 103.665 129.645 ;
        RECT 103.835 128.995 104.095 129.450 ;
        RECT 104.265 129.165 104.565 129.645 ;
        RECT 104.825 129.185 105.385 129.475 ;
        RECT 105.555 129.185 105.805 129.645 ;
        RECT 97.820 128.825 104.565 128.995 ;
        RECT 96.110 128.405 103.230 128.655 ;
        RECT 94.335 127.265 94.505 128.025 ;
        RECT 94.685 127.095 95.015 127.855 ;
        RECT 95.185 127.265 95.455 128.170 ;
        RECT 95.635 127.095 95.930 127.905 ;
        RECT 96.110 127.265 96.355 128.405 ;
        RECT 96.530 127.095 96.790 127.905 ;
        RECT 96.970 127.270 97.220 128.405 ;
        RECT 103.400 128.235 104.565 128.825 ;
        RECT 97.820 128.010 104.565 128.235 ;
        RECT 97.820 127.995 103.225 128.010 ;
        RECT 97.390 127.100 97.650 127.895 ;
        RECT 97.820 127.270 98.080 127.995 ;
        RECT 98.250 127.100 98.510 127.825 ;
        RECT 98.680 127.270 98.940 127.995 ;
        RECT 99.110 127.100 99.370 127.825 ;
        RECT 99.540 127.270 99.800 127.995 ;
        RECT 99.970 127.100 100.230 127.825 ;
        RECT 100.400 127.270 100.660 127.995 ;
        RECT 100.830 127.100 101.075 127.825 ;
        RECT 101.245 127.270 101.505 127.995 ;
        RECT 101.690 127.100 101.935 127.825 ;
        RECT 102.105 127.270 102.365 127.995 ;
        RECT 102.550 127.100 102.795 127.825 ;
        RECT 102.965 127.270 103.225 127.995 ;
        RECT 103.410 127.100 103.665 127.825 ;
        RECT 103.835 127.270 104.125 128.010 ;
        RECT 97.390 127.095 103.665 127.100 ;
        RECT 104.295 127.095 104.565 127.840 ;
        RECT 104.825 127.815 105.075 129.185 ;
        RECT 106.425 129.015 106.755 129.375 ;
        RECT 105.365 128.825 106.755 129.015 ;
        RECT 107.125 129.185 107.685 129.475 ;
        RECT 107.855 129.185 108.105 129.645 ;
        RECT 105.365 128.735 105.535 128.825 ;
        RECT 105.245 128.405 105.535 128.735 ;
        RECT 105.705 128.405 106.045 128.655 ;
        RECT 106.265 128.405 106.940 128.655 ;
        RECT 105.365 128.155 105.535 128.405 ;
        RECT 105.365 127.985 106.305 128.155 ;
        RECT 106.675 128.045 106.940 128.405 ;
        RECT 104.825 127.265 105.285 127.815 ;
        RECT 105.475 127.095 105.805 127.815 ;
        RECT 106.005 127.435 106.305 127.985 ;
        RECT 107.125 127.815 107.375 129.185 ;
        RECT 108.725 129.015 109.055 129.375 ;
        RECT 107.665 128.825 109.055 129.015 ;
        RECT 109.625 129.015 109.955 129.375 ;
        RECT 110.575 129.185 110.825 129.645 ;
        RECT 110.995 129.185 111.555 129.475 ;
        RECT 109.625 128.825 111.015 129.015 ;
        RECT 107.665 128.735 107.835 128.825 ;
        RECT 107.545 128.405 107.835 128.735 ;
        RECT 110.845 128.735 111.015 128.825 ;
        RECT 108.005 128.405 108.345 128.655 ;
        RECT 108.565 128.405 109.240 128.655 ;
        RECT 107.665 128.155 107.835 128.405 ;
        RECT 107.665 127.985 108.605 128.155 ;
        RECT 108.975 128.045 109.240 128.405 ;
        RECT 109.440 128.405 110.115 128.655 ;
        RECT 110.335 128.405 110.675 128.655 ;
        RECT 110.845 128.405 111.135 128.735 ;
        RECT 109.440 128.045 109.705 128.405 ;
        RECT 110.845 128.155 111.015 128.405 ;
        RECT 106.475 127.095 106.755 127.765 ;
        RECT 107.125 127.265 107.585 127.815 ;
        RECT 107.775 127.095 108.105 127.815 ;
        RECT 108.305 127.435 108.605 127.985 ;
        RECT 110.075 127.985 111.015 128.155 ;
        RECT 108.775 127.095 109.055 127.765 ;
        RECT 109.625 127.095 109.905 127.765 ;
        RECT 110.075 127.435 110.375 127.985 ;
        RECT 111.305 127.815 111.555 129.185 ;
        RECT 110.575 127.095 110.905 127.815 ;
        RECT 111.095 127.265 111.555 127.815 ;
        RECT 111.725 129.185 112.285 129.475 ;
        RECT 112.455 129.185 112.705 129.645 ;
        RECT 111.725 127.815 111.975 129.185 ;
        RECT 113.325 129.015 113.655 129.375 ;
        RECT 112.265 128.825 113.655 129.015 ;
        RECT 114.485 128.920 114.775 129.645 ;
        RECT 115.405 128.875 117.995 129.645 ;
        RECT 112.265 128.735 112.435 128.825 ;
        RECT 112.145 128.405 112.435 128.735 ;
        RECT 112.605 128.405 112.945 128.655 ;
        RECT 113.165 128.405 113.840 128.655 ;
        RECT 112.265 128.155 112.435 128.405 ;
        RECT 112.265 127.985 113.205 128.155 ;
        RECT 113.575 128.045 113.840 128.405 ;
        RECT 111.725 127.265 112.185 127.815 ;
        RECT 112.375 127.095 112.705 127.815 ;
        RECT 112.905 127.435 113.205 127.985 ;
        RECT 113.375 127.095 113.655 127.765 ;
        RECT 114.485 127.095 114.775 128.260 ;
        RECT 115.405 128.185 116.615 128.705 ;
        RECT 116.785 128.355 117.995 128.875 ;
        RECT 118.205 128.825 118.435 129.645 ;
        RECT 118.605 128.845 118.935 129.475 ;
        RECT 118.185 128.405 118.515 128.655 ;
        RECT 118.685 128.245 118.935 128.845 ;
        RECT 119.105 128.825 119.315 129.645 ;
        RECT 119.635 129.095 119.805 129.475 ;
        RECT 119.985 129.265 120.315 129.645 ;
        RECT 119.635 128.925 120.300 129.095 ;
        RECT 120.495 128.970 120.755 129.475 ;
        RECT 120.930 129.100 126.275 129.645 ;
        RECT 119.565 128.375 119.895 128.745 ;
        RECT 120.130 128.670 120.300 128.925 ;
        RECT 115.405 127.095 117.995 128.185 ;
        RECT 118.205 127.095 118.435 128.235 ;
        RECT 118.605 127.265 118.935 128.245 ;
        RECT 120.130 128.340 120.415 128.670 ;
        RECT 119.105 127.095 119.315 128.235 ;
        RECT 120.130 128.195 120.300 128.340 ;
        RECT 119.635 128.025 120.300 128.195 ;
        RECT 120.585 128.170 120.755 128.970 ;
        RECT 119.635 127.265 119.805 128.025 ;
        RECT 119.985 127.095 120.315 127.855 ;
        RECT 120.485 127.265 120.755 128.170 ;
        RECT 122.520 127.530 122.870 128.780 ;
        RECT 124.350 128.270 124.690 129.100 ;
        RECT 126.445 128.895 127.655 129.645 ;
        RECT 126.445 128.185 126.965 128.725 ;
        RECT 127.135 128.355 127.655 128.895 ;
        RECT 120.930 127.095 126.275 127.530 ;
        RECT 126.445 127.095 127.655 128.185 ;
        RECT 14.580 126.925 127.740 127.095 ;
        RECT 14.665 125.835 15.875 126.925 ;
        RECT 14.665 125.125 15.185 125.665 ;
        RECT 15.355 125.295 15.875 125.835 ;
        RECT 16.045 125.835 17.255 126.925 ;
        RECT 17.425 125.835 20.935 126.925 ;
        RECT 16.045 125.295 16.565 125.835 ;
        RECT 16.735 125.125 17.255 125.665 ;
        RECT 17.425 125.315 19.115 125.835 ;
        RECT 21.165 125.785 21.375 126.925 ;
        RECT 21.545 125.775 21.875 126.755 ;
        RECT 22.045 125.785 22.275 126.925 ;
        RECT 23.035 125.995 23.205 126.755 ;
        RECT 23.385 126.165 23.715 126.925 ;
        RECT 23.035 125.825 23.700 125.995 ;
        RECT 23.885 125.850 24.155 126.755 ;
        RECT 19.285 125.145 20.935 125.665 ;
        RECT 14.665 124.375 15.875 125.125 ;
        RECT 16.045 124.375 17.255 125.125 ;
        RECT 17.425 124.375 20.935 125.145 ;
        RECT 21.165 124.375 21.375 125.195 ;
        RECT 21.545 125.175 21.795 125.775 ;
        RECT 23.530 125.680 23.700 125.825 ;
        RECT 21.965 125.365 22.295 125.615 ;
        RECT 22.965 125.275 23.295 125.645 ;
        RECT 23.530 125.350 23.815 125.680 ;
        RECT 21.545 124.545 21.875 125.175 ;
        RECT 22.045 124.375 22.275 125.195 ;
        RECT 23.530 125.095 23.700 125.350 ;
        RECT 23.035 124.925 23.700 125.095 ;
        RECT 23.985 125.050 24.155 125.850 ;
        RECT 24.325 125.760 24.615 126.925 ;
        RECT 25.710 126.490 31.055 126.925 ;
        RECT 31.230 126.490 36.575 126.925 ;
        RECT 27.300 125.240 27.650 126.490 ;
        RECT 23.035 124.545 23.205 124.925 ;
        RECT 23.385 124.375 23.715 124.755 ;
        RECT 23.895 124.545 24.155 125.050 ;
        RECT 24.325 124.375 24.615 125.100 ;
        RECT 29.130 124.920 29.470 125.750 ;
        RECT 32.820 125.240 33.170 126.490 ;
        RECT 36.945 126.255 37.225 126.925 ;
        RECT 37.395 126.035 37.695 126.585 ;
        RECT 37.895 126.205 38.225 126.925 ;
        RECT 38.415 126.205 38.875 126.755 ;
        RECT 34.650 124.920 34.990 125.750 ;
        RECT 36.760 125.615 37.025 125.975 ;
        RECT 37.395 125.865 38.335 126.035 ;
        RECT 38.165 125.615 38.335 125.865 ;
        RECT 36.760 125.365 37.435 125.615 ;
        RECT 37.655 125.365 37.995 125.615 ;
        RECT 38.165 125.285 38.455 125.615 ;
        RECT 38.165 125.195 38.335 125.285 ;
        RECT 36.945 125.005 38.335 125.195 ;
        RECT 25.710 124.375 31.055 124.920 ;
        RECT 31.230 124.375 36.575 124.920 ;
        RECT 36.945 124.645 37.275 125.005 ;
        RECT 38.625 124.835 38.875 126.205 ;
        RECT 39.045 125.835 40.255 126.925 ;
        RECT 40.425 126.205 40.885 126.755 ;
        RECT 41.075 126.205 41.405 126.925 ;
        RECT 39.045 125.295 39.565 125.835 ;
        RECT 39.735 125.125 40.255 125.665 ;
        RECT 37.895 124.375 38.145 124.835 ;
        RECT 38.315 124.545 38.875 124.835 ;
        RECT 39.045 124.375 40.255 125.125 ;
        RECT 40.425 124.835 40.675 126.205 ;
        RECT 41.605 126.035 41.905 126.585 ;
        RECT 42.075 126.255 42.355 126.925 ;
        RECT 42.925 126.255 43.205 126.925 ;
        RECT 40.965 125.865 41.905 126.035 ;
        RECT 43.375 126.035 43.675 126.585 ;
        RECT 43.875 126.205 44.205 126.925 ;
        RECT 44.395 126.205 44.855 126.755 ;
        RECT 40.965 125.615 41.135 125.865 ;
        RECT 42.275 125.615 42.540 125.975 ;
        RECT 40.845 125.285 41.135 125.615 ;
        RECT 41.305 125.365 41.645 125.615 ;
        RECT 41.865 125.365 42.540 125.615 ;
        RECT 42.740 125.615 43.005 125.975 ;
        RECT 43.375 125.865 44.315 126.035 ;
        RECT 44.145 125.615 44.315 125.865 ;
        RECT 42.740 125.365 43.415 125.615 ;
        RECT 43.635 125.365 43.975 125.615 ;
        RECT 40.965 125.195 41.135 125.285 ;
        RECT 44.145 125.285 44.435 125.615 ;
        RECT 44.145 125.195 44.315 125.285 ;
        RECT 40.965 125.005 42.355 125.195 ;
        RECT 40.425 124.545 40.985 124.835 ;
        RECT 41.155 124.375 41.405 124.835 ;
        RECT 42.025 124.645 42.355 125.005 ;
        RECT 42.925 125.005 44.315 125.195 ;
        RECT 42.925 124.645 43.255 125.005 ;
        RECT 44.605 124.835 44.855 126.205 ;
        RECT 43.875 124.375 44.125 124.835 ;
        RECT 44.295 124.545 44.855 124.835 ;
        RECT 45.025 126.205 45.485 126.755 ;
        RECT 45.675 126.205 46.005 126.925 ;
        RECT 45.025 124.835 45.275 126.205 ;
        RECT 46.205 126.035 46.505 126.585 ;
        RECT 46.675 126.255 46.955 126.925 ;
        RECT 47.380 126.055 47.665 126.925 ;
        RECT 47.835 126.295 48.095 126.755 ;
        RECT 48.270 126.465 48.525 126.925 ;
        RECT 48.695 126.295 48.955 126.755 ;
        RECT 47.835 126.125 48.955 126.295 ;
        RECT 49.125 126.125 49.435 126.925 ;
        RECT 45.565 125.865 46.505 126.035 ;
        RECT 45.565 125.615 45.735 125.865 ;
        RECT 46.875 125.615 47.140 125.975 ;
        RECT 47.835 125.875 48.095 126.125 ;
        RECT 49.605 125.955 49.915 126.755 ;
        RECT 45.445 125.285 45.735 125.615 ;
        RECT 45.905 125.365 46.245 125.615 ;
        RECT 46.465 125.365 47.140 125.615 ;
        RECT 47.340 125.705 48.095 125.875 ;
        RECT 48.885 125.785 49.915 125.955 ;
        RECT 45.565 125.195 45.735 125.285 ;
        RECT 47.340 125.195 47.745 125.705 ;
        RECT 48.885 125.535 49.055 125.785 ;
        RECT 47.915 125.365 49.055 125.535 ;
        RECT 45.565 125.005 46.955 125.195 ;
        RECT 47.340 125.025 48.990 125.195 ;
        RECT 49.225 125.045 49.575 125.615 ;
        RECT 45.025 124.545 45.585 124.835 ;
        RECT 45.755 124.375 46.005 124.835 ;
        RECT 46.625 124.645 46.955 125.005 ;
        RECT 47.385 124.375 47.665 124.855 ;
        RECT 47.835 124.635 48.095 125.025 ;
        RECT 48.270 124.375 48.525 124.855 ;
        RECT 48.695 124.635 48.990 125.025 ;
        RECT 49.745 124.875 49.915 125.785 ;
        RECT 50.085 125.760 50.375 126.925 ;
        RECT 50.545 125.835 52.215 126.925 ;
        RECT 52.390 126.490 57.735 126.925 ;
        RECT 50.545 125.315 51.295 125.835 ;
        RECT 51.465 125.145 52.215 125.665 ;
        RECT 53.980 125.240 54.330 126.490 ;
        RECT 57.995 125.995 58.165 126.755 ;
        RECT 58.345 126.165 58.675 126.925 ;
        RECT 57.995 125.825 58.660 125.995 ;
        RECT 58.845 125.850 59.115 126.755 ;
        RECT 49.170 124.375 49.445 124.855 ;
        RECT 49.615 124.545 49.915 124.875 ;
        RECT 50.085 124.375 50.375 125.100 ;
        RECT 50.545 124.375 52.215 125.145 ;
        RECT 55.810 124.920 56.150 125.750 ;
        RECT 58.490 125.680 58.660 125.825 ;
        RECT 57.925 125.275 58.255 125.645 ;
        RECT 58.490 125.350 58.775 125.680 ;
        RECT 58.490 125.095 58.660 125.350 ;
        RECT 57.995 124.925 58.660 125.095 ;
        RECT 58.945 125.050 59.115 125.850 ;
        RECT 59.285 126.165 59.800 126.575 ;
        RECT 60.035 126.165 60.205 126.925 ;
        RECT 60.375 126.585 62.405 126.755 ;
        RECT 59.285 125.355 59.625 126.165 ;
        RECT 60.375 125.920 60.545 126.585 ;
        RECT 60.940 126.245 62.065 126.415 ;
        RECT 59.795 125.730 60.545 125.920 ;
        RECT 60.715 125.905 61.725 126.075 ;
        RECT 59.285 125.185 60.515 125.355 ;
        RECT 52.390 124.375 57.735 124.920 ;
        RECT 57.995 124.545 58.165 124.925 ;
        RECT 58.345 124.375 58.675 124.755 ;
        RECT 58.855 124.545 59.115 125.050 ;
        RECT 59.560 124.580 59.805 125.185 ;
        RECT 60.025 124.375 60.535 124.910 ;
        RECT 60.715 124.545 60.905 125.905 ;
        RECT 61.075 125.565 61.350 125.705 ;
        RECT 61.075 125.395 61.355 125.565 ;
        RECT 61.075 124.545 61.350 125.395 ;
        RECT 61.555 125.105 61.725 125.905 ;
        RECT 61.895 125.115 62.065 126.245 ;
        RECT 62.235 125.615 62.405 126.585 ;
        RECT 62.575 125.785 62.745 126.925 ;
        RECT 62.915 125.785 63.250 126.755 ;
        RECT 62.235 125.285 62.430 125.615 ;
        RECT 62.655 125.285 62.910 125.615 ;
        RECT 62.655 125.115 62.825 125.285 ;
        RECT 63.080 125.115 63.250 125.785 ;
        RECT 63.425 125.835 64.635 126.925 ;
        RECT 64.805 125.835 68.315 126.925 ;
        RECT 63.425 125.295 63.945 125.835 ;
        RECT 64.115 125.125 64.635 125.665 ;
        RECT 64.805 125.315 66.495 125.835 ;
        RECT 68.545 125.785 68.755 126.925 ;
        RECT 68.925 125.775 69.255 126.755 ;
        RECT 69.425 125.785 69.655 126.925 ;
        RECT 70.415 125.995 70.585 126.755 ;
        RECT 70.765 126.165 71.095 126.925 ;
        RECT 70.415 125.825 71.080 125.995 ;
        RECT 71.265 125.850 71.535 126.755 ;
        RECT 66.665 125.145 68.315 125.665 ;
        RECT 61.895 124.945 62.825 125.115 ;
        RECT 61.895 124.910 62.070 124.945 ;
        RECT 61.540 124.545 62.070 124.910 ;
        RECT 62.495 124.375 62.825 124.775 ;
        RECT 62.995 124.545 63.250 125.115 ;
        RECT 63.425 124.375 64.635 125.125 ;
        RECT 64.805 124.375 68.315 125.145 ;
        RECT 68.545 124.375 68.755 125.195 ;
        RECT 68.925 125.175 69.175 125.775 ;
        RECT 70.910 125.680 71.080 125.825 ;
        RECT 69.345 125.365 69.675 125.615 ;
        RECT 70.345 125.275 70.675 125.645 ;
        RECT 70.910 125.350 71.195 125.680 ;
        RECT 68.925 124.545 69.255 125.175 ;
        RECT 69.425 124.375 69.655 125.195 ;
        RECT 70.910 125.095 71.080 125.350 ;
        RECT 70.415 124.925 71.080 125.095 ;
        RECT 71.365 125.050 71.535 125.850 ;
        RECT 70.415 124.545 70.585 124.925 ;
        RECT 70.765 124.375 71.095 124.755 ;
        RECT 71.275 124.545 71.535 125.050 ;
        RECT 72.625 125.955 72.935 126.755 ;
        RECT 73.105 126.125 73.415 126.925 ;
        RECT 73.585 126.295 73.845 126.755 ;
        RECT 74.015 126.465 74.270 126.925 ;
        RECT 74.445 126.295 74.705 126.755 ;
        RECT 73.585 126.125 74.705 126.295 ;
        RECT 72.625 125.785 73.655 125.955 ;
        RECT 72.625 124.875 72.795 125.785 ;
        RECT 72.965 125.045 73.315 125.615 ;
        RECT 73.485 125.535 73.655 125.785 ;
        RECT 74.445 125.875 74.705 126.125 ;
        RECT 74.875 126.055 75.160 126.925 ;
        RECT 74.445 125.705 75.200 125.875 ;
        RECT 75.845 125.760 76.135 126.925 ;
        RECT 76.305 125.835 77.975 126.925 ;
        RECT 78.520 126.585 78.775 126.615 ;
        RECT 78.435 126.415 78.775 126.585 ;
        RECT 78.520 125.945 78.775 126.415 ;
        RECT 78.955 126.125 79.240 126.925 ;
        RECT 79.420 126.205 79.750 126.715 ;
        RECT 73.485 125.365 74.625 125.535 ;
        RECT 74.795 125.195 75.200 125.705 ;
        RECT 76.305 125.315 77.055 125.835 ;
        RECT 73.550 125.025 75.200 125.195 ;
        RECT 77.225 125.145 77.975 125.665 ;
        RECT 72.625 124.545 72.925 124.875 ;
        RECT 73.095 124.375 73.370 124.855 ;
        RECT 73.550 124.635 73.845 125.025 ;
        RECT 74.015 124.375 74.270 124.855 ;
        RECT 74.445 124.635 74.705 125.025 ;
        RECT 74.875 124.375 75.155 124.855 ;
        RECT 75.845 124.375 76.135 125.100 ;
        RECT 76.305 124.375 77.975 125.145 ;
        RECT 78.520 125.085 78.700 125.945 ;
        RECT 79.420 125.615 79.670 126.205 ;
        RECT 80.020 126.055 80.190 126.665 ;
        RECT 80.360 126.235 80.690 126.925 ;
        RECT 80.920 126.375 81.160 126.665 ;
        RECT 81.360 126.545 81.780 126.925 ;
        RECT 81.960 126.455 82.590 126.705 ;
        RECT 83.060 126.545 83.390 126.925 ;
        RECT 81.960 126.375 82.130 126.455 ;
        RECT 83.560 126.375 83.730 126.665 ;
        RECT 83.910 126.545 84.290 126.925 ;
        RECT 84.530 126.540 85.360 126.710 ;
        RECT 80.920 126.205 82.130 126.375 ;
        RECT 78.870 125.285 79.670 125.615 ;
        RECT 78.520 124.555 78.775 125.085 ;
        RECT 78.955 124.375 79.240 124.835 ;
        RECT 79.420 124.635 79.670 125.285 ;
        RECT 79.870 126.035 80.190 126.055 ;
        RECT 79.870 125.865 81.790 126.035 ;
        RECT 79.870 124.970 80.060 125.865 ;
        RECT 81.960 125.695 82.130 126.205 ;
        RECT 82.300 125.945 82.820 126.255 ;
        RECT 80.230 125.525 82.130 125.695 ;
        RECT 80.230 125.465 80.560 125.525 ;
        RECT 80.710 125.295 81.040 125.355 ;
        RECT 80.380 125.025 81.040 125.295 ;
        RECT 79.870 124.640 80.190 124.970 ;
        RECT 80.370 124.375 81.030 124.855 ;
        RECT 81.230 124.765 81.400 125.525 ;
        RECT 82.300 125.355 82.480 125.765 ;
        RECT 81.570 125.185 81.900 125.305 ;
        RECT 82.650 125.185 82.820 125.945 ;
        RECT 81.570 125.015 82.820 125.185 ;
        RECT 82.990 126.125 84.360 126.375 ;
        RECT 82.990 125.355 83.180 126.125 ;
        RECT 84.110 125.865 84.360 126.125 ;
        RECT 83.350 125.695 83.600 125.855 ;
        RECT 84.530 125.695 84.700 126.540 ;
        RECT 85.595 126.255 85.765 126.755 ;
        RECT 85.935 126.425 86.265 126.925 ;
        RECT 84.870 125.865 85.370 126.245 ;
        RECT 85.595 126.085 86.290 126.255 ;
        RECT 83.350 125.525 84.700 125.695 ;
        RECT 84.280 125.485 84.700 125.525 ;
        RECT 82.990 125.015 83.410 125.355 ;
        RECT 83.700 125.025 84.110 125.355 ;
        RECT 81.230 124.595 82.080 124.765 ;
        RECT 82.640 124.375 82.960 124.835 ;
        RECT 83.160 124.585 83.410 125.015 ;
        RECT 83.700 124.375 84.110 124.815 ;
        RECT 84.280 124.755 84.450 125.485 ;
        RECT 84.620 124.935 84.970 125.305 ;
        RECT 85.150 124.995 85.370 125.865 ;
        RECT 85.540 125.295 85.950 125.915 ;
        RECT 86.120 125.115 86.290 126.085 ;
        RECT 85.595 124.925 86.290 125.115 ;
        RECT 84.280 124.555 85.295 124.755 ;
        RECT 85.595 124.595 85.765 124.925 ;
        RECT 85.935 124.375 86.265 124.755 ;
        RECT 86.480 124.635 86.705 126.755 ;
        RECT 86.875 126.425 87.205 126.925 ;
        RECT 87.375 126.255 87.545 126.755 ;
        RECT 86.880 126.085 87.545 126.255 ;
        RECT 86.880 125.095 87.110 126.085 ;
        RECT 87.280 125.265 87.630 125.915 ;
        RECT 87.805 125.835 89.475 126.925 ;
        RECT 89.735 126.255 89.905 126.755 ;
        RECT 90.075 126.425 90.405 126.925 ;
        RECT 89.735 126.085 90.400 126.255 ;
        RECT 87.805 125.315 88.555 125.835 ;
        RECT 88.725 125.145 89.475 125.665 ;
        RECT 89.650 125.265 90.000 125.915 ;
        RECT 86.880 124.925 87.545 125.095 ;
        RECT 86.875 124.375 87.205 124.755 ;
        RECT 87.375 124.635 87.545 124.925 ;
        RECT 87.805 124.375 89.475 125.145 ;
        RECT 90.170 125.095 90.400 126.085 ;
        RECT 89.735 124.925 90.400 125.095 ;
        RECT 89.735 124.635 89.905 124.925 ;
        RECT 90.075 124.375 90.405 124.755 ;
        RECT 90.575 124.635 90.800 126.755 ;
        RECT 91.015 126.425 91.345 126.925 ;
        RECT 91.515 126.255 91.685 126.755 ;
        RECT 91.920 126.540 92.750 126.710 ;
        RECT 92.990 126.545 93.370 126.925 ;
        RECT 90.990 126.085 91.685 126.255 ;
        RECT 90.990 125.115 91.160 126.085 ;
        RECT 91.330 125.295 91.740 125.915 ;
        RECT 91.910 125.865 92.410 126.245 ;
        RECT 90.990 124.925 91.685 125.115 ;
        RECT 91.910 124.995 92.130 125.865 ;
        RECT 92.580 125.695 92.750 126.540 ;
        RECT 93.550 126.375 93.720 126.665 ;
        RECT 93.890 126.545 94.220 126.925 ;
        RECT 94.690 126.455 95.320 126.705 ;
        RECT 95.500 126.545 95.920 126.925 ;
        RECT 95.150 126.375 95.320 126.455 ;
        RECT 96.120 126.375 96.360 126.665 ;
        RECT 92.920 126.125 94.290 126.375 ;
        RECT 92.920 125.865 93.170 126.125 ;
        RECT 93.680 125.695 93.930 125.855 ;
        RECT 92.580 125.525 93.930 125.695 ;
        RECT 92.580 125.485 93.000 125.525 ;
        RECT 92.310 124.935 92.660 125.305 ;
        RECT 91.015 124.375 91.345 124.755 ;
        RECT 91.515 124.595 91.685 124.925 ;
        RECT 92.830 124.755 93.000 125.485 ;
        RECT 94.100 125.355 94.290 126.125 ;
        RECT 93.170 125.025 93.580 125.355 ;
        RECT 93.870 125.015 94.290 125.355 ;
        RECT 94.460 125.945 94.980 126.255 ;
        RECT 95.150 126.205 96.360 126.375 ;
        RECT 96.590 126.235 96.920 126.925 ;
        RECT 94.460 125.185 94.630 125.945 ;
        RECT 94.800 125.355 94.980 125.765 ;
        RECT 95.150 125.695 95.320 126.205 ;
        RECT 97.090 126.055 97.260 126.665 ;
        RECT 97.530 126.205 97.860 126.715 ;
        RECT 97.090 126.035 97.410 126.055 ;
        RECT 95.490 125.865 97.410 126.035 ;
        RECT 95.150 125.525 97.050 125.695 ;
        RECT 95.380 125.185 95.710 125.305 ;
        RECT 94.460 125.015 95.710 125.185 ;
        RECT 91.985 124.555 93.000 124.755 ;
        RECT 93.170 124.375 93.580 124.815 ;
        RECT 93.870 124.585 94.120 125.015 ;
        RECT 94.320 124.375 94.640 124.835 ;
        RECT 95.880 124.765 96.050 125.525 ;
        RECT 96.720 125.465 97.050 125.525 ;
        RECT 96.240 125.295 96.570 125.355 ;
        RECT 96.240 125.025 96.900 125.295 ;
        RECT 97.220 124.970 97.410 125.865 ;
        RECT 95.200 124.595 96.050 124.765 ;
        RECT 96.250 124.375 96.910 124.855 ;
        RECT 97.090 124.640 97.410 124.970 ;
        RECT 97.610 125.615 97.860 126.205 ;
        RECT 98.040 126.125 98.325 126.925 ;
        RECT 98.505 126.585 98.760 126.615 ;
        RECT 98.505 126.415 98.845 126.585 ;
        RECT 98.505 125.945 98.760 126.415 ;
        RECT 99.505 126.255 99.785 126.925 ;
        RECT 99.955 126.035 100.255 126.585 ;
        RECT 100.455 126.205 100.785 126.925 ;
        RECT 100.975 126.205 101.435 126.755 ;
        RECT 97.610 125.285 98.410 125.615 ;
        RECT 97.610 124.635 97.860 125.285 ;
        RECT 98.580 125.085 98.760 125.945 ;
        RECT 99.320 125.615 99.585 125.975 ;
        RECT 99.955 125.865 100.895 126.035 ;
        RECT 100.725 125.615 100.895 125.865 ;
        RECT 99.320 125.365 99.995 125.615 ;
        RECT 100.215 125.365 100.555 125.615 ;
        RECT 100.725 125.285 101.015 125.615 ;
        RECT 100.725 125.195 100.895 125.285 ;
        RECT 98.040 124.375 98.325 124.835 ;
        RECT 98.505 124.555 98.760 125.085 ;
        RECT 99.505 125.005 100.895 125.195 ;
        RECT 99.505 124.645 99.835 125.005 ;
        RECT 101.185 124.835 101.435 126.205 ;
        RECT 101.605 125.760 101.895 126.925 ;
        RECT 102.065 125.835 105.575 126.925 ;
        RECT 105.750 126.490 111.095 126.925 ;
        RECT 102.065 125.315 103.755 125.835 ;
        RECT 103.925 125.145 105.575 125.665 ;
        RECT 107.340 125.240 107.690 126.490 ;
        RECT 111.265 126.165 111.780 126.575 ;
        RECT 112.015 126.165 112.185 126.925 ;
        RECT 112.355 126.585 114.385 126.755 ;
        RECT 100.455 124.375 100.705 124.835 ;
        RECT 100.875 124.545 101.435 124.835 ;
        RECT 101.605 124.375 101.895 125.100 ;
        RECT 102.065 124.375 105.575 125.145 ;
        RECT 109.170 124.920 109.510 125.750 ;
        RECT 111.265 125.355 111.605 126.165 ;
        RECT 112.355 125.920 112.525 126.585 ;
        RECT 112.920 126.245 114.045 126.415 ;
        RECT 111.775 125.730 112.525 125.920 ;
        RECT 112.695 125.905 113.705 126.075 ;
        RECT 111.265 125.185 112.495 125.355 ;
        RECT 105.750 124.375 111.095 124.920 ;
        RECT 111.540 124.580 111.785 125.185 ;
        RECT 112.005 124.375 112.515 124.910 ;
        RECT 112.695 124.545 112.885 125.905 ;
        RECT 113.055 124.885 113.330 125.705 ;
        RECT 113.535 125.105 113.705 125.905 ;
        RECT 113.875 125.115 114.045 126.245 ;
        RECT 114.215 125.615 114.385 126.585 ;
        RECT 114.555 125.785 114.725 126.925 ;
        RECT 114.895 125.785 115.230 126.755 ;
        RECT 114.215 125.285 114.410 125.615 ;
        RECT 114.635 125.285 114.890 125.615 ;
        RECT 114.635 125.115 114.805 125.285 ;
        RECT 115.060 125.115 115.230 125.785 ;
        RECT 113.875 124.945 114.805 125.115 ;
        RECT 113.875 124.910 114.050 124.945 ;
        RECT 113.055 124.715 113.335 124.885 ;
        RECT 113.055 124.545 113.330 124.715 ;
        RECT 113.520 124.545 114.050 124.910 ;
        RECT 114.475 124.375 114.805 124.775 ;
        RECT 114.975 124.545 115.230 125.115 ;
        RECT 115.780 125.945 116.035 126.615 ;
        RECT 116.215 126.125 116.500 126.925 ;
        RECT 116.680 126.205 117.010 126.715 ;
        RECT 115.780 125.085 115.960 125.945 ;
        RECT 116.680 125.615 116.930 126.205 ;
        RECT 117.280 126.055 117.450 126.665 ;
        RECT 117.620 126.235 117.950 126.925 ;
        RECT 118.180 126.375 118.420 126.665 ;
        RECT 118.620 126.545 119.040 126.925 ;
        RECT 119.220 126.455 119.850 126.705 ;
        RECT 120.320 126.545 120.650 126.925 ;
        RECT 119.220 126.375 119.390 126.455 ;
        RECT 120.820 126.375 120.990 126.665 ;
        RECT 121.170 126.545 121.550 126.925 ;
        RECT 121.790 126.540 122.620 126.710 ;
        RECT 118.180 126.205 119.390 126.375 ;
        RECT 116.130 125.285 116.930 125.615 ;
        RECT 115.780 124.885 116.035 125.085 ;
        RECT 115.695 124.715 116.035 124.885 ;
        RECT 115.780 124.555 116.035 124.715 ;
        RECT 116.215 124.375 116.500 124.835 ;
        RECT 116.680 124.635 116.930 125.285 ;
        RECT 117.130 126.035 117.450 126.055 ;
        RECT 117.130 125.865 119.050 126.035 ;
        RECT 117.130 124.970 117.320 125.865 ;
        RECT 119.220 125.695 119.390 126.205 ;
        RECT 119.560 125.945 120.080 126.255 ;
        RECT 117.490 125.525 119.390 125.695 ;
        RECT 117.490 125.465 117.820 125.525 ;
        RECT 117.970 125.295 118.300 125.355 ;
        RECT 117.640 125.025 118.300 125.295 ;
        RECT 117.130 124.640 117.450 124.970 ;
        RECT 117.630 124.375 118.290 124.855 ;
        RECT 118.490 124.765 118.660 125.525 ;
        RECT 119.560 125.355 119.740 125.765 ;
        RECT 118.830 125.185 119.160 125.305 ;
        RECT 119.910 125.185 120.080 125.945 ;
        RECT 118.830 125.015 120.080 125.185 ;
        RECT 120.250 126.125 121.620 126.375 ;
        RECT 120.250 125.355 120.440 126.125 ;
        RECT 121.370 125.865 121.620 126.125 ;
        RECT 120.610 125.695 120.860 125.855 ;
        RECT 121.790 125.695 121.960 126.540 ;
        RECT 122.855 126.255 123.025 126.755 ;
        RECT 123.195 126.425 123.525 126.925 ;
        RECT 122.130 125.865 122.630 126.245 ;
        RECT 122.855 126.085 123.550 126.255 ;
        RECT 120.610 125.525 121.960 125.695 ;
        RECT 121.540 125.485 121.960 125.525 ;
        RECT 120.250 125.015 120.670 125.355 ;
        RECT 120.960 125.025 121.370 125.355 ;
        RECT 118.490 124.595 119.340 124.765 ;
        RECT 119.900 124.375 120.220 124.835 ;
        RECT 120.420 124.585 120.670 125.015 ;
        RECT 120.960 124.375 121.370 124.815 ;
        RECT 121.540 124.755 121.710 125.485 ;
        RECT 121.880 124.935 122.230 125.305 ;
        RECT 122.410 124.995 122.630 125.865 ;
        RECT 122.800 125.295 123.210 125.915 ;
        RECT 123.380 125.115 123.550 126.085 ;
        RECT 122.855 124.925 123.550 125.115 ;
        RECT 121.540 124.555 122.555 124.755 ;
        RECT 122.855 124.595 123.025 124.925 ;
        RECT 123.195 124.375 123.525 124.755 ;
        RECT 123.740 124.635 123.965 126.755 ;
        RECT 124.135 126.425 124.465 126.925 ;
        RECT 124.635 126.255 124.805 126.755 ;
        RECT 124.140 126.085 124.805 126.255 ;
        RECT 124.140 125.095 124.370 126.085 ;
        RECT 124.540 125.265 124.890 125.915 ;
        RECT 125.065 125.835 126.275 126.925 ;
        RECT 126.445 125.835 127.655 126.925 ;
        RECT 125.065 125.295 125.585 125.835 ;
        RECT 125.755 125.125 126.275 125.665 ;
        RECT 126.445 125.295 126.965 125.835 ;
        RECT 127.135 125.125 127.655 125.665 ;
        RECT 124.140 124.925 124.805 125.095 ;
        RECT 124.135 124.375 124.465 124.755 ;
        RECT 124.635 124.635 124.805 124.925 ;
        RECT 125.065 124.375 126.275 125.125 ;
        RECT 126.445 124.375 127.655 125.125 ;
        RECT 14.580 124.205 127.740 124.375 ;
        RECT 14.665 123.455 15.875 124.205 ;
        RECT 16.045 123.455 17.255 124.205 ;
        RECT 17.430 123.660 22.775 124.205 ;
        RECT 14.665 122.915 15.185 123.455 ;
        RECT 15.355 122.745 15.875 123.285 ;
        RECT 14.665 121.655 15.875 122.745 ;
        RECT 16.045 122.745 16.565 123.285 ;
        RECT 16.735 122.915 17.255 123.455 ;
        RECT 16.045 121.655 17.255 122.745 ;
        RECT 19.020 122.090 19.370 123.340 ;
        RECT 20.850 122.830 21.190 123.660 ;
        RECT 23.220 123.395 23.465 124.000 ;
        RECT 23.685 123.670 24.195 124.205 ;
        RECT 22.945 123.225 24.175 123.395 ;
        RECT 22.945 122.415 23.285 123.225 ;
        RECT 23.455 122.660 24.205 122.850 ;
        RECT 17.430 121.655 22.775 122.090 ;
        RECT 22.945 122.005 23.460 122.415 ;
        RECT 23.695 121.655 23.865 122.415 ;
        RECT 24.035 121.995 24.205 122.660 ;
        RECT 24.375 122.675 24.565 124.035 ;
        RECT 24.735 123.865 25.010 124.035 ;
        RECT 24.735 123.695 25.015 123.865 ;
        RECT 24.735 122.875 25.010 123.695 ;
        RECT 25.200 123.670 25.730 124.035 ;
        RECT 26.155 123.805 26.485 124.205 ;
        RECT 25.555 123.635 25.730 123.670 ;
        RECT 25.215 122.675 25.385 123.475 ;
        RECT 24.375 122.505 25.385 122.675 ;
        RECT 25.555 123.465 26.485 123.635 ;
        RECT 26.655 123.465 26.910 124.035 ;
        RECT 27.550 123.660 32.895 124.205 ;
        RECT 25.555 122.335 25.725 123.465 ;
        RECT 26.315 123.295 26.485 123.465 ;
        RECT 24.600 122.165 25.725 122.335 ;
        RECT 25.895 122.965 26.090 123.295 ;
        RECT 26.315 122.965 26.570 123.295 ;
        RECT 25.895 121.995 26.065 122.965 ;
        RECT 26.740 122.795 26.910 123.465 ;
        RECT 24.035 121.825 26.065 121.995 ;
        RECT 26.235 121.655 26.405 122.795 ;
        RECT 26.575 121.825 26.910 122.795 ;
        RECT 29.140 122.090 29.490 123.340 ;
        RECT 30.970 122.830 31.310 123.660 ;
        RECT 33.340 123.395 33.585 124.000 ;
        RECT 33.805 123.670 34.315 124.205 ;
        RECT 33.065 123.225 34.295 123.395 ;
        RECT 33.065 122.415 33.405 123.225 ;
        RECT 33.575 122.660 34.325 122.850 ;
        RECT 27.550 121.655 32.895 122.090 ;
        RECT 33.065 122.005 33.580 122.415 ;
        RECT 33.815 121.655 33.985 122.415 ;
        RECT 34.155 121.995 34.325 122.660 ;
        RECT 34.495 122.675 34.685 124.035 ;
        RECT 34.855 123.185 35.130 124.035 ;
        RECT 35.320 123.670 35.850 124.035 ;
        RECT 36.275 123.805 36.605 124.205 ;
        RECT 35.675 123.635 35.850 123.670 ;
        RECT 34.855 123.015 35.135 123.185 ;
        RECT 34.855 122.875 35.130 123.015 ;
        RECT 35.335 122.675 35.505 123.475 ;
        RECT 34.495 122.505 35.505 122.675 ;
        RECT 35.675 123.465 36.605 123.635 ;
        RECT 36.775 123.465 37.030 124.035 ;
        RECT 37.205 123.480 37.495 124.205 ;
        RECT 35.675 122.335 35.845 123.465 ;
        RECT 36.435 123.295 36.605 123.465 ;
        RECT 34.720 122.165 35.845 122.335 ;
        RECT 36.015 122.965 36.210 123.295 ;
        RECT 36.435 122.965 36.690 123.295 ;
        RECT 36.015 121.995 36.185 122.965 ;
        RECT 36.860 122.795 37.030 123.465 ;
        RECT 38.125 123.435 41.635 124.205 ;
        RECT 41.810 123.660 47.155 124.205 ;
        RECT 47.330 123.660 52.675 124.205 ;
        RECT 53.220 123.865 53.475 124.025 ;
        RECT 53.135 123.695 53.475 123.865 ;
        RECT 53.655 123.745 53.940 124.205 ;
        RECT 34.155 121.825 36.185 121.995 ;
        RECT 36.355 121.655 36.525 122.795 ;
        RECT 36.695 121.825 37.030 122.795 ;
        RECT 37.205 121.655 37.495 122.820 ;
        RECT 38.125 122.745 39.815 123.265 ;
        RECT 39.985 122.915 41.635 123.435 ;
        RECT 38.125 121.655 41.635 122.745 ;
        RECT 43.400 122.090 43.750 123.340 ;
        RECT 45.230 122.830 45.570 123.660 ;
        RECT 48.920 122.090 49.270 123.340 ;
        RECT 50.750 122.830 51.090 123.660 ;
        RECT 53.220 123.495 53.475 123.695 ;
        RECT 53.220 122.635 53.400 123.495 ;
        RECT 54.120 123.295 54.370 123.945 ;
        RECT 53.570 122.965 54.370 123.295 ;
        RECT 41.810 121.655 47.155 122.090 ;
        RECT 47.330 121.655 52.675 122.090 ;
        RECT 53.220 121.965 53.475 122.635 ;
        RECT 53.655 121.655 53.940 122.455 ;
        RECT 54.120 122.375 54.370 122.965 ;
        RECT 54.570 123.610 54.890 123.940 ;
        RECT 55.070 123.725 55.730 124.205 ;
        RECT 55.930 123.815 56.780 123.985 ;
        RECT 54.570 122.715 54.760 123.610 ;
        RECT 55.080 123.285 55.740 123.555 ;
        RECT 55.410 123.225 55.740 123.285 ;
        RECT 54.930 123.055 55.260 123.115 ;
        RECT 55.930 123.055 56.100 123.815 ;
        RECT 57.340 123.745 57.660 124.205 ;
        RECT 57.860 123.565 58.110 123.995 ;
        RECT 58.400 123.765 58.810 124.205 ;
        RECT 58.980 123.825 59.995 124.025 ;
        RECT 56.270 123.395 57.520 123.565 ;
        RECT 56.270 123.275 56.600 123.395 ;
        RECT 54.930 122.885 56.830 123.055 ;
        RECT 54.570 122.545 56.490 122.715 ;
        RECT 54.570 122.525 54.890 122.545 ;
        RECT 54.120 121.865 54.450 122.375 ;
        RECT 54.720 121.915 54.890 122.525 ;
        RECT 56.660 122.375 56.830 122.885 ;
        RECT 57.000 122.815 57.180 123.225 ;
        RECT 57.350 122.635 57.520 123.395 ;
        RECT 55.060 121.655 55.390 122.345 ;
        RECT 55.620 122.205 56.830 122.375 ;
        RECT 57.000 122.325 57.520 122.635 ;
        RECT 57.690 123.225 58.110 123.565 ;
        RECT 58.400 123.225 58.810 123.555 ;
        RECT 57.690 122.455 57.880 123.225 ;
        RECT 58.980 123.095 59.150 123.825 ;
        RECT 60.295 123.655 60.465 123.985 ;
        RECT 60.635 123.825 60.965 124.205 ;
        RECT 59.320 123.275 59.670 123.645 ;
        RECT 58.980 123.055 59.400 123.095 ;
        RECT 58.050 122.885 59.400 123.055 ;
        RECT 58.050 122.725 58.300 122.885 ;
        RECT 58.810 122.455 59.060 122.715 ;
        RECT 57.690 122.205 59.060 122.455 ;
        RECT 55.620 121.915 55.860 122.205 ;
        RECT 56.660 122.125 56.830 122.205 ;
        RECT 56.060 121.655 56.480 122.035 ;
        RECT 56.660 121.875 57.290 122.125 ;
        RECT 57.760 121.655 58.090 122.035 ;
        RECT 58.260 121.915 58.430 122.205 ;
        RECT 59.230 122.040 59.400 122.885 ;
        RECT 59.850 122.715 60.070 123.585 ;
        RECT 60.295 123.465 60.990 123.655 ;
        RECT 59.570 122.335 60.070 122.715 ;
        RECT 60.240 122.665 60.650 123.285 ;
        RECT 60.820 122.495 60.990 123.465 ;
        RECT 60.295 122.325 60.990 122.495 ;
        RECT 58.610 121.655 58.990 122.035 ;
        RECT 59.230 121.870 60.060 122.040 ;
        RECT 60.295 121.825 60.465 122.325 ;
        RECT 60.635 121.655 60.965 122.155 ;
        RECT 61.180 121.825 61.405 123.945 ;
        RECT 61.575 123.825 61.905 124.205 ;
        RECT 62.075 123.655 62.245 123.945 ;
        RECT 61.580 123.485 62.245 123.655 ;
        RECT 61.580 122.495 61.810 123.485 ;
        RECT 62.965 123.480 63.255 124.205 ;
        RECT 64.160 123.395 64.405 124.000 ;
        RECT 64.625 123.670 65.135 124.205 ;
        RECT 61.980 122.665 62.330 123.315 ;
        RECT 63.885 123.225 65.115 123.395 ;
        RECT 61.580 122.325 62.245 122.495 ;
        RECT 61.575 121.655 61.905 122.155 ;
        RECT 62.075 121.825 62.245 122.325 ;
        RECT 62.965 121.655 63.255 122.820 ;
        RECT 63.885 122.415 64.225 123.225 ;
        RECT 64.395 122.660 65.145 122.850 ;
        RECT 63.885 122.005 64.400 122.415 ;
        RECT 64.635 121.655 64.805 122.415 ;
        RECT 64.975 121.995 65.145 122.660 ;
        RECT 65.315 122.675 65.505 124.035 ;
        RECT 65.675 123.865 65.950 124.035 ;
        RECT 65.675 123.695 65.955 123.865 ;
        RECT 65.675 122.875 65.950 123.695 ;
        RECT 66.140 123.670 66.670 124.035 ;
        RECT 67.095 123.805 67.425 124.205 ;
        RECT 66.495 123.635 66.670 123.670 ;
        RECT 66.155 122.675 66.325 123.475 ;
        RECT 65.315 122.505 66.325 122.675 ;
        RECT 66.495 123.465 67.425 123.635 ;
        RECT 67.595 123.465 67.850 124.035 ;
        RECT 66.495 122.335 66.665 123.465 ;
        RECT 67.255 123.295 67.425 123.465 ;
        RECT 65.540 122.165 66.665 122.335 ;
        RECT 66.835 122.965 67.030 123.295 ;
        RECT 67.255 122.965 67.510 123.295 ;
        RECT 66.835 121.995 67.005 122.965 ;
        RECT 67.680 122.795 67.850 123.465 ;
        RECT 68.025 123.435 70.615 124.205 ;
        RECT 70.790 123.660 76.135 124.205 ;
        RECT 76.310 123.660 81.655 124.205 ;
        RECT 64.975 121.825 67.005 121.995 ;
        RECT 67.175 121.655 67.345 122.795 ;
        RECT 67.515 121.825 67.850 122.795 ;
        RECT 68.025 122.745 69.235 123.265 ;
        RECT 69.405 122.915 70.615 123.435 ;
        RECT 68.025 121.655 70.615 122.745 ;
        RECT 72.380 122.090 72.730 123.340 ;
        RECT 74.210 122.830 74.550 123.660 ;
        RECT 77.900 122.090 78.250 123.340 ;
        RECT 79.730 122.830 80.070 123.660 ;
        RECT 81.885 123.385 82.095 124.205 ;
        RECT 82.265 123.405 82.595 124.035 ;
        RECT 82.265 122.805 82.515 123.405 ;
        RECT 82.765 123.385 82.995 124.205 ;
        RECT 83.755 123.655 83.925 124.035 ;
        RECT 84.105 123.825 84.435 124.205 ;
        RECT 83.755 123.485 84.420 123.655 ;
        RECT 84.615 123.530 84.875 124.035 ;
        RECT 82.685 122.965 83.015 123.215 ;
        RECT 83.685 122.935 84.015 123.305 ;
        RECT 84.250 123.230 84.420 123.485 ;
        RECT 84.250 122.900 84.535 123.230 ;
        RECT 70.790 121.655 76.135 122.090 ;
        RECT 76.310 121.655 81.655 122.090 ;
        RECT 81.885 121.655 82.095 122.795 ;
        RECT 82.265 121.825 82.595 122.805 ;
        RECT 82.765 121.655 82.995 122.795 ;
        RECT 84.250 122.755 84.420 122.900 ;
        RECT 83.755 122.585 84.420 122.755 ;
        RECT 84.705 122.730 84.875 123.530 ;
        RECT 85.045 123.435 88.555 124.205 ;
        RECT 88.725 123.480 89.015 124.205 ;
        RECT 89.185 123.435 92.695 124.205 ;
        RECT 83.755 121.825 83.925 122.585 ;
        RECT 84.105 121.655 84.435 122.415 ;
        RECT 84.605 121.825 84.875 122.730 ;
        RECT 85.045 122.745 86.735 123.265 ;
        RECT 86.905 122.915 88.555 123.435 ;
        RECT 85.045 121.655 88.555 122.745 ;
        RECT 88.725 121.655 89.015 122.820 ;
        RECT 89.185 122.745 90.875 123.265 ;
        RECT 91.045 122.915 92.695 123.435 ;
        RECT 92.905 123.385 93.135 124.205 ;
        RECT 93.305 123.405 93.635 124.035 ;
        RECT 92.885 122.965 93.215 123.215 ;
        RECT 93.385 122.805 93.635 123.405 ;
        RECT 93.805 123.385 94.015 124.205 ;
        RECT 94.245 123.455 95.455 124.205 ;
        RECT 89.185 121.655 92.695 122.745 ;
        RECT 92.905 121.655 93.135 122.795 ;
        RECT 93.305 121.825 93.635 122.805 ;
        RECT 93.805 121.655 94.015 122.795 ;
        RECT 94.245 122.745 94.765 123.285 ;
        RECT 94.935 122.915 95.455 123.455 ;
        RECT 95.625 123.435 99.135 124.205 ;
        RECT 99.310 123.660 104.655 124.205 ;
        RECT 104.830 123.660 110.175 124.205 ;
        RECT 95.625 122.745 97.315 123.265 ;
        RECT 97.485 122.915 99.135 123.435 ;
        RECT 94.245 121.655 95.455 122.745 ;
        RECT 95.625 121.655 99.135 122.745 ;
        RECT 100.900 122.090 101.250 123.340 ;
        RECT 102.730 122.830 103.070 123.660 ;
        RECT 106.420 122.090 106.770 123.340 ;
        RECT 108.250 122.830 108.590 123.660 ;
        RECT 110.620 123.395 110.865 124.000 ;
        RECT 111.085 123.670 111.595 124.205 ;
        RECT 110.345 123.225 111.575 123.395 ;
        RECT 110.345 122.415 110.685 123.225 ;
        RECT 110.855 122.660 111.605 122.850 ;
        RECT 99.310 121.655 104.655 122.090 ;
        RECT 104.830 121.655 110.175 122.090 ;
        RECT 110.345 122.005 110.860 122.415 ;
        RECT 111.095 121.655 111.265 122.415 ;
        RECT 111.435 121.995 111.605 122.660 ;
        RECT 111.775 122.675 111.965 124.035 ;
        RECT 112.135 123.185 112.410 124.035 ;
        RECT 112.600 123.670 113.130 124.035 ;
        RECT 113.555 123.805 113.885 124.205 ;
        RECT 112.955 123.635 113.130 123.670 ;
        RECT 112.135 123.015 112.415 123.185 ;
        RECT 112.135 122.875 112.410 123.015 ;
        RECT 112.615 122.675 112.785 123.475 ;
        RECT 111.775 122.505 112.785 122.675 ;
        RECT 112.955 123.465 113.885 123.635 ;
        RECT 114.055 123.465 114.310 124.035 ;
        RECT 114.485 123.480 114.775 124.205 ;
        RECT 115.780 123.495 116.035 124.025 ;
        RECT 116.215 123.745 116.500 124.205 ;
        RECT 112.955 122.335 113.125 123.465 ;
        RECT 113.715 123.295 113.885 123.465 ;
        RECT 112.000 122.165 113.125 122.335 ;
        RECT 113.295 122.965 113.490 123.295 ;
        RECT 113.715 122.965 113.970 123.295 ;
        RECT 113.295 121.995 113.465 122.965 ;
        RECT 114.140 122.795 114.310 123.465 ;
        RECT 115.780 123.185 115.960 123.495 ;
        RECT 116.680 123.295 116.930 123.945 ;
        RECT 115.695 123.015 115.960 123.185 ;
        RECT 111.435 121.825 113.465 121.995 ;
        RECT 113.635 121.655 113.805 122.795 ;
        RECT 113.975 121.825 114.310 122.795 ;
        RECT 114.485 121.655 114.775 122.820 ;
        RECT 115.780 122.635 115.960 123.015 ;
        RECT 116.130 122.965 116.930 123.295 ;
        RECT 115.780 121.965 116.035 122.635 ;
        RECT 116.215 121.655 116.500 122.455 ;
        RECT 116.680 122.375 116.930 122.965 ;
        RECT 117.130 123.610 117.450 123.940 ;
        RECT 117.630 123.725 118.290 124.205 ;
        RECT 118.490 123.815 119.340 123.985 ;
        RECT 117.130 122.715 117.320 123.610 ;
        RECT 117.640 123.285 118.300 123.555 ;
        RECT 117.970 123.225 118.300 123.285 ;
        RECT 117.490 123.055 117.820 123.115 ;
        RECT 118.490 123.055 118.660 123.815 ;
        RECT 119.900 123.745 120.220 124.205 ;
        RECT 120.420 123.565 120.670 123.995 ;
        RECT 120.960 123.765 121.370 124.205 ;
        RECT 121.540 123.825 122.555 124.025 ;
        RECT 118.830 123.395 120.080 123.565 ;
        RECT 118.830 123.275 119.160 123.395 ;
        RECT 117.490 122.885 119.390 123.055 ;
        RECT 117.130 122.545 119.050 122.715 ;
        RECT 117.130 122.525 117.450 122.545 ;
        RECT 116.680 121.865 117.010 122.375 ;
        RECT 117.280 121.915 117.450 122.525 ;
        RECT 119.220 122.375 119.390 122.885 ;
        RECT 119.560 122.815 119.740 123.225 ;
        RECT 119.910 122.635 120.080 123.395 ;
        RECT 117.620 121.655 117.950 122.345 ;
        RECT 118.180 122.205 119.390 122.375 ;
        RECT 119.560 122.325 120.080 122.635 ;
        RECT 120.250 123.225 120.670 123.565 ;
        RECT 120.960 123.225 121.370 123.555 ;
        RECT 120.250 122.455 120.440 123.225 ;
        RECT 121.540 123.095 121.710 123.825 ;
        RECT 122.855 123.655 123.025 123.985 ;
        RECT 123.195 123.825 123.525 124.205 ;
        RECT 121.880 123.275 122.230 123.645 ;
        RECT 121.540 123.055 121.960 123.095 ;
        RECT 120.610 122.885 121.960 123.055 ;
        RECT 120.610 122.725 120.860 122.885 ;
        RECT 121.370 122.455 121.620 122.715 ;
        RECT 120.250 122.205 121.620 122.455 ;
        RECT 118.180 121.915 118.420 122.205 ;
        RECT 119.220 122.125 119.390 122.205 ;
        RECT 118.620 121.655 119.040 122.035 ;
        RECT 119.220 121.875 119.850 122.125 ;
        RECT 120.320 121.655 120.650 122.035 ;
        RECT 120.820 121.915 120.990 122.205 ;
        RECT 121.790 122.040 121.960 122.885 ;
        RECT 122.410 122.715 122.630 123.585 ;
        RECT 122.855 123.465 123.550 123.655 ;
        RECT 122.130 122.335 122.630 122.715 ;
        RECT 122.800 122.665 123.210 123.285 ;
        RECT 123.380 122.495 123.550 123.465 ;
        RECT 122.855 122.325 123.550 122.495 ;
        RECT 121.170 121.655 121.550 122.035 ;
        RECT 121.790 121.870 122.620 122.040 ;
        RECT 122.855 121.825 123.025 122.325 ;
        RECT 123.195 121.655 123.525 122.155 ;
        RECT 123.740 121.825 123.965 123.945 ;
        RECT 124.135 123.825 124.465 124.205 ;
        RECT 124.635 123.655 124.805 123.945 ;
        RECT 124.140 123.485 124.805 123.655 ;
        RECT 124.140 122.495 124.370 123.485 ;
        RECT 125.065 123.455 126.275 124.205 ;
        RECT 126.445 123.455 127.655 124.205 ;
        RECT 124.540 122.665 124.890 123.315 ;
        RECT 125.065 122.745 125.585 123.285 ;
        RECT 125.755 122.915 126.275 123.455 ;
        RECT 126.445 122.745 126.965 123.285 ;
        RECT 127.135 122.915 127.655 123.455 ;
        RECT 124.140 122.325 124.805 122.495 ;
        RECT 124.135 121.655 124.465 122.155 ;
        RECT 124.635 121.825 124.805 122.325 ;
        RECT 125.065 121.655 126.275 122.745 ;
        RECT 126.445 121.655 127.655 122.745 ;
        RECT 14.580 121.485 127.740 121.655 ;
        RECT 14.665 120.395 15.875 121.485 ;
        RECT 14.665 119.685 15.185 120.225 ;
        RECT 15.355 119.855 15.875 120.395 ;
        RECT 16.505 120.395 20.015 121.485 ;
        RECT 16.505 119.875 18.195 120.395 ;
        RECT 20.190 120.345 20.525 121.315 ;
        RECT 20.695 120.345 20.865 121.485 ;
        RECT 21.035 121.145 23.065 121.315 ;
        RECT 18.365 119.705 20.015 120.225 ;
        RECT 14.665 118.935 15.875 119.685 ;
        RECT 16.505 118.935 20.015 119.705 ;
        RECT 20.190 119.675 20.360 120.345 ;
        RECT 21.035 120.175 21.205 121.145 ;
        RECT 20.530 119.845 20.785 120.175 ;
        RECT 21.010 119.845 21.205 120.175 ;
        RECT 21.375 120.805 22.500 120.975 ;
        RECT 20.615 119.675 20.785 119.845 ;
        RECT 21.375 119.675 21.545 120.805 ;
        RECT 20.190 119.105 20.445 119.675 ;
        RECT 20.615 119.505 21.545 119.675 ;
        RECT 21.715 120.465 22.725 120.635 ;
        RECT 21.715 119.665 21.885 120.465 ;
        RECT 22.090 119.785 22.365 120.265 ;
        RECT 22.085 119.615 22.365 119.785 ;
        RECT 21.370 119.470 21.545 119.505 ;
        RECT 20.615 118.935 20.945 119.335 ;
        RECT 21.370 119.105 21.900 119.470 ;
        RECT 22.090 119.105 22.365 119.615 ;
        RECT 22.535 119.105 22.725 120.465 ;
        RECT 22.895 120.480 23.065 121.145 ;
        RECT 23.235 120.725 23.405 121.485 ;
        RECT 23.640 120.725 24.155 121.135 ;
        RECT 22.895 120.290 23.645 120.480 ;
        RECT 23.815 119.915 24.155 120.725 ;
        RECT 24.325 120.320 24.615 121.485 ;
        RECT 24.785 120.395 25.995 121.485 ;
        RECT 26.165 120.410 26.435 121.315 ;
        RECT 26.605 120.725 26.935 121.485 ;
        RECT 27.115 120.555 27.285 121.315 ;
        RECT 22.925 119.745 24.155 119.915 ;
        RECT 24.785 119.855 25.305 120.395 ;
        RECT 22.905 118.935 23.415 119.470 ;
        RECT 23.635 119.140 23.880 119.745 ;
        RECT 25.475 119.685 25.995 120.225 ;
        RECT 24.325 118.935 24.615 119.660 ;
        RECT 24.785 118.935 25.995 119.685 ;
        RECT 26.165 119.610 26.335 120.410 ;
        RECT 26.620 120.385 27.285 120.555 ;
        RECT 27.545 120.395 30.135 121.485 ;
        RECT 30.680 121.145 30.935 121.175 ;
        RECT 30.595 120.975 30.935 121.145 ;
        RECT 30.680 120.505 30.935 120.975 ;
        RECT 31.115 120.685 31.400 121.485 ;
        RECT 31.580 120.765 31.910 121.275 ;
        RECT 26.620 120.240 26.790 120.385 ;
        RECT 26.505 119.910 26.790 120.240 ;
        RECT 26.620 119.655 26.790 119.910 ;
        RECT 27.025 119.835 27.355 120.205 ;
        RECT 27.545 119.875 28.755 120.395 ;
        RECT 28.925 119.705 30.135 120.225 ;
        RECT 26.165 119.105 26.425 119.610 ;
        RECT 26.620 119.485 27.285 119.655 ;
        RECT 26.605 118.935 26.935 119.315 ;
        RECT 27.115 119.105 27.285 119.485 ;
        RECT 27.545 118.935 30.135 119.705 ;
        RECT 30.680 119.645 30.860 120.505 ;
        RECT 31.580 120.175 31.830 120.765 ;
        RECT 32.180 120.615 32.350 121.225 ;
        RECT 32.520 120.795 32.850 121.485 ;
        RECT 33.080 120.935 33.320 121.225 ;
        RECT 33.520 121.105 33.940 121.485 ;
        RECT 34.120 121.015 34.750 121.265 ;
        RECT 35.220 121.105 35.550 121.485 ;
        RECT 34.120 120.935 34.290 121.015 ;
        RECT 35.720 120.935 35.890 121.225 ;
        RECT 36.070 121.105 36.450 121.485 ;
        RECT 36.690 121.100 37.520 121.270 ;
        RECT 33.080 120.765 34.290 120.935 ;
        RECT 31.030 119.845 31.830 120.175 ;
        RECT 30.680 119.115 30.935 119.645 ;
        RECT 31.115 118.935 31.400 119.395 ;
        RECT 31.580 119.195 31.830 119.845 ;
        RECT 32.030 120.595 32.350 120.615 ;
        RECT 32.030 120.425 33.950 120.595 ;
        RECT 32.030 119.530 32.220 120.425 ;
        RECT 34.120 120.255 34.290 120.765 ;
        RECT 34.460 120.505 34.980 120.815 ;
        RECT 32.390 120.085 34.290 120.255 ;
        RECT 32.390 120.025 32.720 120.085 ;
        RECT 32.870 119.855 33.200 119.915 ;
        RECT 32.540 119.585 33.200 119.855 ;
        RECT 32.030 119.200 32.350 119.530 ;
        RECT 32.530 118.935 33.190 119.415 ;
        RECT 33.390 119.325 33.560 120.085 ;
        RECT 34.460 119.915 34.640 120.325 ;
        RECT 33.730 119.745 34.060 119.865 ;
        RECT 34.810 119.745 34.980 120.505 ;
        RECT 33.730 119.575 34.980 119.745 ;
        RECT 35.150 120.685 36.520 120.935 ;
        RECT 35.150 119.915 35.340 120.685 ;
        RECT 36.270 120.425 36.520 120.685 ;
        RECT 35.510 120.255 35.760 120.415 ;
        RECT 36.690 120.255 36.860 121.100 ;
        RECT 37.755 120.815 37.925 121.315 ;
        RECT 38.095 120.985 38.425 121.485 ;
        RECT 37.030 120.425 37.530 120.805 ;
        RECT 37.755 120.645 38.450 120.815 ;
        RECT 35.510 120.085 36.860 120.255 ;
        RECT 36.440 120.045 36.860 120.085 ;
        RECT 35.150 119.575 35.570 119.915 ;
        RECT 35.860 119.585 36.270 119.915 ;
        RECT 33.390 119.155 34.240 119.325 ;
        RECT 34.800 118.935 35.120 119.395 ;
        RECT 35.320 119.145 35.570 119.575 ;
        RECT 35.860 118.935 36.270 119.375 ;
        RECT 36.440 119.315 36.610 120.045 ;
        RECT 36.780 119.495 37.130 119.865 ;
        RECT 37.310 119.555 37.530 120.425 ;
        RECT 37.700 119.855 38.110 120.475 ;
        RECT 38.280 119.675 38.450 120.645 ;
        RECT 37.755 119.485 38.450 119.675 ;
        RECT 36.440 119.115 37.455 119.315 ;
        RECT 37.755 119.155 37.925 119.485 ;
        RECT 38.095 118.935 38.425 119.315 ;
        RECT 38.640 119.195 38.865 121.315 ;
        RECT 39.035 120.985 39.365 121.485 ;
        RECT 39.535 120.815 39.705 121.315 ;
        RECT 39.040 120.645 39.705 120.815 ;
        RECT 39.040 119.655 39.270 120.645 ;
        RECT 39.440 119.825 39.790 120.475 ;
        RECT 39.970 120.345 40.305 121.315 ;
        RECT 40.475 120.345 40.645 121.485 ;
        RECT 40.815 121.145 42.845 121.315 ;
        RECT 39.970 119.675 40.140 120.345 ;
        RECT 40.815 120.175 40.985 121.145 ;
        RECT 40.310 119.845 40.565 120.175 ;
        RECT 40.790 119.845 40.985 120.175 ;
        RECT 41.155 120.805 42.280 120.975 ;
        RECT 40.395 119.675 40.565 119.845 ;
        RECT 41.155 119.675 41.325 120.805 ;
        RECT 39.040 119.485 39.705 119.655 ;
        RECT 39.035 118.935 39.365 119.315 ;
        RECT 39.535 119.195 39.705 119.485 ;
        RECT 39.970 119.105 40.225 119.675 ;
        RECT 40.395 119.505 41.325 119.675 ;
        RECT 41.495 120.465 42.505 120.635 ;
        RECT 41.495 119.665 41.665 120.465 ;
        RECT 41.870 120.125 42.145 120.265 ;
        RECT 41.865 119.955 42.145 120.125 ;
        RECT 41.150 119.470 41.325 119.505 ;
        RECT 40.395 118.935 40.725 119.335 ;
        RECT 41.150 119.105 41.680 119.470 ;
        RECT 41.870 119.105 42.145 119.955 ;
        RECT 42.315 119.105 42.505 120.465 ;
        RECT 42.675 120.480 42.845 121.145 ;
        RECT 43.015 120.725 43.185 121.485 ;
        RECT 43.420 120.725 43.935 121.135 ;
        RECT 42.675 120.290 43.425 120.480 ;
        RECT 43.595 119.915 43.935 120.725 ;
        RECT 42.705 119.745 43.935 119.915 ;
        RECT 44.565 120.410 44.835 121.315 ;
        RECT 45.005 120.725 45.335 121.485 ;
        RECT 45.515 120.555 45.685 121.315 ;
        RECT 42.685 118.935 43.195 119.470 ;
        RECT 43.415 119.140 43.660 119.745 ;
        RECT 44.565 119.610 44.735 120.410 ;
        RECT 45.020 120.385 45.685 120.555 ;
        RECT 45.945 120.725 46.460 121.135 ;
        RECT 46.695 120.725 46.865 121.485 ;
        RECT 47.035 121.145 49.065 121.315 ;
        RECT 45.020 120.240 45.190 120.385 ;
        RECT 44.905 119.910 45.190 120.240 ;
        RECT 45.020 119.655 45.190 119.910 ;
        RECT 45.425 119.835 45.755 120.205 ;
        RECT 45.945 119.915 46.285 120.725 ;
        RECT 47.035 120.480 47.205 121.145 ;
        RECT 47.600 120.805 48.725 120.975 ;
        RECT 46.455 120.290 47.205 120.480 ;
        RECT 47.375 120.465 48.385 120.635 ;
        RECT 45.945 119.745 47.175 119.915 ;
        RECT 44.565 119.105 44.825 119.610 ;
        RECT 45.020 119.485 45.685 119.655 ;
        RECT 45.005 118.935 45.335 119.315 ;
        RECT 45.515 119.105 45.685 119.485 ;
        RECT 46.220 119.140 46.465 119.745 ;
        RECT 46.685 118.935 47.195 119.470 ;
        RECT 47.375 119.105 47.565 120.465 ;
        RECT 47.735 120.125 48.010 120.265 ;
        RECT 47.735 119.955 48.015 120.125 ;
        RECT 47.735 119.105 48.010 119.955 ;
        RECT 48.215 119.665 48.385 120.465 ;
        RECT 48.555 119.675 48.725 120.805 ;
        RECT 48.895 120.175 49.065 121.145 ;
        RECT 49.235 120.345 49.405 121.485 ;
        RECT 49.575 120.345 49.910 121.315 ;
        RECT 48.895 119.845 49.090 120.175 ;
        RECT 49.315 119.845 49.570 120.175 ;
        RECT 49.315 119.675 49.485 119.845 ;
        RECT 49.740 119.675 49.910 120.345 ;
        RECT 50.085 120.320 50.375 121.485 ;
        RECT 50.585 120.345 50.815 121.485 ;
        RECT 50.985 120.335 51.315 121.315 ;
        RECT 51.485 120.345 51.695 121.485 ;
        RECT 51.925 120.395 53.135 121.485 ;
        RECT 50.565 119.925 50.895 120.175 ;
        RECT 48.555 119.505 49.485 119.675 ;
        RECT 48.555 119.470 48.730 119.505 ;
        RECT 48.200 119.105 48.730 119.470 ;
        RECT 49.155 118.935 49.485 119.335 ;
        RECT 49.655 119.105 49.910 119.675 ;
        RECT 50.085 118.935 50.375 119.660 ;
        RECT 50.585 118.935 50.815 119.755 ;
        RECT 51.065 119.735 51.315 120.335 ;
        RECT 51.925 119.855 52.445 120.395 ;
        RECT 53.455 120.335 53.785 121.485 ;
        RECT 53.955 120.465 54.125 121.315 ;
        RECT 54.295 120.685 54.625 121.485 ;
        RECT 54.795 120.465 54.965 121.315 ;
        RECT 55.145 120.685 55.385 121.485 ;
        RECT 55.555 120.505 55.885 121.315 ;
        RECT 53.955 120.295 54.965 120.465 ;
        RECT 55.170 120.335 55.885 120.505 ;
        RECT 57.045 120.345 57.255 121.485 ;
        RECT 57.425 120.335 57.755 121.315 ;
        RECT 57.925 120.345 58.155 121.485 ;
        RECT 59.660 121.145 59.915 121.175 ;
        RECT 59.575 120.975 59.915 121.145 ;
        RECT 59.660 120.505 59.915 120.975 ;
        RECT 60.095 120.685 60.380 121.485 ;
        RECT 60.560 120.765 60.890 121.275 ;
        RECT 50.985 119.105 51.315 119.735 ;
        RECT 51.485 118.935 51.695 119.755 ;
        RECT 52.615 119.685 53.135 120.225 ;
        RECT 53.955 120.125 54.450 120.295 ;
        RECT 53.955 119.955 54.455 120.125 ;
        RECT 55.170 120.095 55.340 120.335 ;
        RECT 53.955 119.755 54.450 119.955 ;
        RECT 54.840 119.925 55.340 120.095 ;
        RECT 55.510 119.925 55.890 120.165 ;
        RECT 55.170 119.755 55.340 119.925 ;
        RECT 51.925 118.935 53.135 119.685 ;
        RECT 53.455 118.935 53.785 119.735 ;
        RECT 53.955 119.585 54.965 119.755 ;
        RECT 55.170 119.585 55.805 119.755 ;
        RECT 53.955 119.105 54.125 119.585 ;
        RECT 54.295 118.935 54.625 119.415 ;
        RECT 54.795 119.105 54.965 119.585 ;
        RECT 55.215 118.935 55.455 119.415 ;
        RECT 55.635 119.105 55.805 119.585 ;
        RECT 57.045 118.935 57.255 119.755 ;
        RECT 57.425 119.735 57.675 120.335 ;
        RECT 57.845 119.925 58.175 120.175 ;
        RECT 57.425 119.105 57.755 119.735 ;
        RECT 57.925 118.935 58.155 119.755 ;
        RECT 59.660 119.645 59.840 120.505 ;
        RECT 60.560 120.175 60.810 120.765 ;
        RECT 61.160 120.615 61.330 121.225 ;
        RECT 61.500 120.795 61.830 121.485 ;
        RECT 62.060 120.935 62.300 121.225 ;
        RECT 62.500 121.105 62.920 121.485 ;
        RECT 63.100 121.015 63.730 121.265 ;
        RECT 64.200 121.105 64.530 121.485 ;
        RECT 63.100 120.935 63.270 121.015 ;
        RECT 64.700 120.935 64.870 121.225 ;
        RECT 65.050 121.105 65.430 121.485 ;
        RECT 65.670 121.100 66.500 121.270 ;
        RECT 62.060 120.765 63.270 120.935 ;
        RECT 60.010 119.845 60.810 120.175 ;
        RECT 59.660 119.115 59.915 119.645 ;
        RECT 60.095 118.935 60.380 119.395 ;
        RECT 60.560 119.195 60.810 119.845 ;
        RECT 61.010 120.595 61.330 120.615 ;
        RECT 61.010 120.425 62.930 120.595 ;
        RECT 61.010 119.530 61.200 120.425 ;
        RECT 63.100 120.255 63.270 120.765 ;
        RECT 63.440 120.505 63.960 120.815 ;
        RECT 61.370 120.085 63.270 120.255 ;
        RECT 61.370 120.025 61.700 120.085 ;
        RECT 61.850 119.855 62.180 119.915 ;
        RECT 61.520 119.585 62.180 119.855 ;
        RECT 61.010 119.200 61.330 119.530 ;
        RECT 61.510 118.935 62.170 119.415 ;
        RECT 62.370 119.325 62.540 120.085 ;
        RECT 63.440 119.915 63.620 120.325 ;
        RECT 62.710 119.745 63.040 119.865 ;
        RECT 63.790 119.745 63.960 120.505 ;
        RECT 62.710 119.575 63.960 119.745 ;
        RECT 64.130 120.685 65.500 120.935 ;
        RECT 64.130 119.915 64.320 120.685 ;
        RECT 65.250 120.425 65.500 120.685 ;
        RECT 64.490 120.255 64.740 120.415 ;
        RECT 65.670 120.255 65.840 121.100 ;
        RECT 66.735 120.815 66.905 121.315 ;
        RECT 67.075 120.985 67.405 121.485 ;
        RECT 66.010 120.425 66.510 120.805 ;
        RECT 66.735 120.645 67.430 120.815 ;
        RECT 64.490 120.085 65.840 120.255 ;
        RECT 65.420 120.045 65.840 120.085 ;
        RECT 64.130 119.575 64.550 119.915 ;
        RECT 64.840 119.585 65.250 119.915 ;
        RECT 62.370 119.155 63.220 119.325 ;
        RECT 63.780 118.935 64.100 119.395 ;
        RECT 64.300 119.145 64.550 119.575 ;
        RECT 64.840 118.935 65.250 119.375 ;
        RECT 65.420 119.315 65.590 120.045 ;
        RECT 65.760 119.495 66.110 119.865 ;
        RECT 66.290 119.555 66.510 120.425 ;
        RECT 66.680 119.855 67.090 120.475 ;
        RECT 67.260 119.675 67.430 120.645 ;
        RECT 66.735 119.485 67.430 119.675 ;
        RECT 65.420 119.115 66.435 119.315 ;
        RECT 66.735 119.155 66.905 119.485 ;
        RECT 67.075 118.935 67.405 119.315 ;
        RECT 67.620 119.195 67.845 121.315 ;
        RECT 68.015 120.985 68.345 121.485 ;
        RECT 68.515 120.815 68.685 121.315 ;
        RECT 68.020 120.645 68.685 120.815 ;
        RECT 68.020 119.655 68.250 120.645 ;
        RECT 68.420 119.825 68.770 120.475 ;
        RECT 68.945 120.410 69.215 121.315 ;
        RECT 69.385 120.725 69.715 121.485 ;
        RECT 69.895 120.555 70.065 121.315 ;
        RECT 68.020 119.485 68.685 119.655 ;
        RECT 68.015 118.935 68.345 119.315 ;
        RECT 68.515 119.195 68.685 119.485 ;
        RECT 68.945 119.610 69.115 120.410 ;
        RECT 69.400 120.385 70.065 120.555 ;
        RECT 70.785 120.395 74.295 121.485 ;
        RECT 69.400 120.240 69.570 120.385 ;
        RECT 69.285 119.910 69.570 120.240 ;
        RECT 69.400 119.655 69.570 119.910 ;
        RECT 69.805 119.835 70.135 120.205 ;
        RECT 70.785 119.875 72.475 120.395 ;
        RECT 74.505 120.345 74.735 121.485 ;
        RECT 74.905 120.335 75.235 121.315 ;
        RECT 75.405 120.345 75.615 121.485 ;
        RECT 72.645 119.705 74.295 120.225 ;
        RECT 74.485 119.925 74.815 120.175 ;
        RECT 68.945 119.105 69.205 119.610 ;
        RECT 69.400 119.485 70.065 119.655 ;
        RECT 69.385 118.935 69.715 119.315 ;
        RECT 69.895 119.105 70.065 119.485 ;
        RECT 70.785 118.935 74.295 119.705 ;
        RECT 74.505 118.935 74.735 119.755 ;
        RECT 74.985 119.735 75.235 120.335 ;
        RECT 75.845 120.320 76.135 121.485 ;
        RECT 76.765 120.725 77.280 121.135 ;
        RECT 77.515 120.725 77.685 121.485 ;
        RECT 77.855 121.145 79.885 121.315 ;
        RECT 76.765 119.915 77.105 120.725 ;
        RECT 77.855 120.480 78.025 121.145 ;
        RECT 78.420 120.805 79.545 120.975 ;
        RECT 77.275 120.290 78.025 120.480 ;
        RECT 78.195 120.465 79.205 120.635 ;
        RECT 74.905 119.105 75.235 119.735 ;
        RECT 75.405 118.935 75.615 119.755 ;
        RECT 76.765 119.745 77.995 119.915 ;
        RECT 75.845 118.935 76.135 119.660 ;
        RECT 77.040 119.140 77.285 119.745 ;
        RECT 77.505 118.935 78.015 119.470 ;
        RECT 78.195 119.105 78.385 120.465 ;
        RECT 78.555 119.445 78.830 120.265 ;
        RECT 79.035 119.665 79.205 120.465 ;
        RECT 79.375 119.675 79.545 120.805 ;
        RECT 79.715 120.175 79.885 121.145 ;
        RECT 80.055 120.345 80.225 121.485 ;
        RECT 80.395 120.345 80.730 121.315 ;
        RECT 79.715 119.845 79.910 120.175 ;
        RECT 80.135 119.845 80.390 120.175 ;
        RECT 80.135 119.675 80.305 119.845 ;
        RECT 80.560 119.675 80.730 120.345 ;
        RECT 79.375 119.505 80.305 119.675 ;
        RECT 79.375 119.470 79.550 119.505 ;
        RECT 78.555 119.275 78.835 119.445 ;
        RECT 78.555 119.105 78.830 119.275 ;
        RECT 79.020 119.105 79.550 119.470 ;
        RECT 79.975 118.935 80.305 119.335 ;
        RECT 80.475 119.105 80.730 119.675 ;
        RECT 80.905 120.410 81.175 121.315 ;
        RECT 81.345 120.725 81.675 121.485 ;
        RECT 81.855 120.555 82.025 121.315 ;
        RECT 80.905 119.610 81.075 120.410 ;
        RECT 81.360 120.385 82.025 120.555 ;
        RECT 81.360 120.240 81.530 120.385 ;
        RECT 82.345 120.345 82.555 121.485 ;
        RECT 81.245 119.910 81.530 120.240 ;
        RECT 82.725 120.335 83.055 121.315 ;
        RECT 83.225 120.345 83.455 121.485 ;
        RECT 84.215 120.555 84.385 121.315 ;
        RECT 84.565 120.725 84.895 121.485 ;
        RECT 84.215 120.385 84.880 120.555 ;
        RECT 85.065 120.410 85.335 121.315 ;
        RECT 85.510 121.050 90.855 121.485 ;
        RECT 81.360 119.655 81.530 119.910 ;
        RECT 81.765 119.835 82.095 120.205 ;
        RECT 80.905 119.105 81.165 119.610 ;
        RECT 81.360 119.485 82.025 119.655 ;
        RECT 81.345 118.935 81.675 119.315 ;
        RECT 81.855 119.105 82.025 119.485 ;
        RECT 82.345 118.935 82.555 119.755 ;
        RECT 82.725 119.735 82.975 120.335 ;
        RECT 84.710 120.240 84.880 120.385 ;
        RECT 83.145 119.925 83.475 120.175 ;
        RECT 84.145 119.835 84.475 120.205 ;
        RECT 84.710 119.910 84.995 120.240 ;
        RECT 82.725 119.105 83.055 119.735 ;
        RECT 83.225 118.935 83.455 119.755 ;
        RECT 84.710 119.655 84.880 119.910 ;
        RECT 84.215 119.485 84.880 119.655 ;
        RECT 85.165 119.610 85.335 120.410 ;
        RECT 87.100 119.800 87.450 121.050 ;
        RECT 91.030 120.345 91.365 121.315 ;
        RECT 91.535 120.345 91.705 121.485 ;
        RECT 91.875 121.145 93.905 121.315 ;
        RECT 84.215 119.105 84.385 119.485 ;
        RECT 84.565 118.935 84.895 119.315 ;
        RECT 85.075 119.105 85.335 119.610 ;
        RECT 88.930 119.480 89.270 120.310 ;
        RECT 91.030 119.675 91.200 120.345 ;
        RECT 91.875 120.175 92.045 121.145 ;
        RECT 91.370 119.845 91.625 120.175 ;
        RECT 91.850 119.845 92.045 120.175 ;
        RECT 92.215 120.805 93.340 120.975 ;
        RECT 91.455 119.675 91.625 119.845 ;
        RECT 92.215 119.675 92.385 120.805 ;
        RECT 85.510 118.935 90.855 119.480 ;
        RECT 91.030 119.105 91.285 119.675 ;
        RECT 91.455 119.505 92.385 119.675 ;
        RECT 92.555 120.465 93.565 120.635 ;
        RECT 92.555 119.665 92.725 120.465 ;
        RECT 92.210 119.470 92.385 119.505 ;
        RECT 91.455 118.935 91.785 119.335 ;
        RECT 92.210 119.105 92.740 119.470 ;
        RECT 92.930 119.445 93.205 120.265 ;
        RECT 92.925 119.275 93.205 119.445 ;
        RECT 92.930 119.105 93.205 119.275 ;
        RECT 93.375 119.105 93.565 120.465 ;
        RECT 93.735 120.480 93.905 121.145 ;
        RECT 94.075 120.725 94.245 121.485 ;
        RECT 94.480 120.725 94.995 121.135 ;
        RECT 93.735 120.290 94.485 120.480 ;
        RECT 94.655 119.915 94.995 120.725 ;
        RECT 93.765 119.745 94.995 119.915 ;
        RECT 95.625 120.395 97.295 121.485 ;
        RECT 97.465 120.725 97.980 121.135 ;
        RECT 98.215 120.725 98.385 121.485 ;
        RECT 98.555 121.145 100.585 121.315 ;
        RECT 95.625 119.875 96.375 120.395 ;
        RECT 93.745 118.935 94.255 119.470 ;
        RECT 94.475 119.140 94.720 119.745 ;
        RECT 96.545 119.705 97.295 120.225 ;
        RECT 97.465 119.915 97.805 120.725 ;
        RECT 98.555 120.480 98.725 121.145 ;
        RECT 99.120 120.805 100.245 120.975 ;
        RECT 97.975 120.290 98.725 120.480 ;
        RECT 98.895 120.465 99.905 120.635 ;
        RECT 97.465 119.745 98.695 119.915 ;
        RECT 95.625 118.935 97.295 119.705 ;
        RECT 97.740 119.140 97.985 119.745 ;
        RECT 98.205 118.935 98.715 119.470 ;
        RECT 98.895 119.105 99.085 120.465 ;
        RECT 99.255 120.125 99.530 120.265 ;
        RECT 99.255 119.955 99.535 120.125 ;
        RECT 99.255 119.105 99.530 119.955 ;
        RECT 99.735 119.665 99.905 120.465 ;
        RECT 100.075 119.675 100.245 120.805 ;
        RECT 100.415 120.175 100.585 121.145 ;
        RECT 100.755 120.345 100.925 121.485 ;
        RECT 101.095 120.345 101.430 121.315 ;
        RECT 100.415 119.845 100.610 120.175 ;
        RECT 100.835 119.845 101.090 120.175 ;
        RECT 100.835 119.675 101.005 119.845 ;
        RECT 101.260 119.675 101.430 120.345 ;
        RECT 101.605 120.320 101.895 121.485 ;
        RECT 102.065 120.395 103.275 121.485 ;
        RECT 102.065 119.855 102.585 120.395 ;
        RECT 103.485 120.345 103.715 121.485 ;
        RECT 103.885 120.335 104.215 121.315 ;
        RECT 104.385 120.345 104.595 121.485 ;
        RECT 104.825 120.725 105.340 121.135 ;
        RECT 105.575 120.725 105.745 121.485 ;
        RECT 105.915 121.145 107.945 121.315 ;
        RECT 102.755 119.685 103.275 120.225 ;
        RECT 103.465 119.925 103.795 120.175 ;
        RECT 100.075 119.505 101.005 119.675 ;
        RECT 100.075 119.470 100.250 119.505 ;
        RECT 99.720 119.105 100.250 119.470 ;
        RECT 100.675 118.935 101.005 119.335 ;
        RECT 101.175 119.105 101.430 119.675 ;
        RECT 101.605 118.935 101.895 119.660 ;
        RECT 102.065 118.935 103.275 119.685 ;
        RECT 103.485 118.935 103.715 119.755 ;
        RECT 103.965 119.735 104.215 120.335 ;
        RECT 104.825 119.915 105.165 120.725 ;
        RECT 105.915 120.480 106.085 121.145 ;
        RECT 106.480 120.805 107.605 120.975 ;
        RECT 105.335 120.290 106.085 120.480 ;
        RECT 106.255 120.465 107.265 120.635 ;
        RECT 103.885 119.105 104.215 119.735 ;
        RECT 104.385 118.935 104.595 119.755 ;
        RECT 104.825 119.745 106.055 119.915 ;
        RECT 105.100 119.140 105.345 119.745 ;
        RECT 105.565 118.935 106.075 119.470 ;
        RECT 106.255 119.105 106.445 120.465 ;
        RECT 106.615 119.785 106.890 120.265 ;
        RECT 106.615 119.615 106.895 119.785 ;
        RECT 107.095 119.665 107.265 120.465 ;
        RECT 107.435 119.675 107.605 120.805 ;
        RECT 107.775 120.175 107.945 121.145 ;
        RECT 108.115 120.345 108.285 121.485 ;
        RECT 108.455 120.345 108.790 121.315 ;
        RECT 109.340 120.505 109.595 121.175 ;
        RECT 109.775 120.685 110.060 121.485 ;
        RECT 110.240 120.765 110.570 121.275 ;
        RECT 109.340 120.465 109.520 120.505 ;
        RECT 107.775 119.845 107.970 120.175 ;
        RECT 108.195 119.845 108.450 120.175 ;
        RECT 108.195 119.675 108.365 119.845 ;
        RECT 108.620 119.675 108.790 120.345 ;
        RECT 109.255 120.295 109.520 120.465 ;
        RECT 106.615 119.105 106.890 119.615 ;
        RECT 107.435 119.505 108.365 119.675 ;
        RECT 107.435 119.470 107.610 119.505 ;
        RECT 107.080 119.105 107.610 119.470 ;
        RECT 108.035 118.935 108.365 119.335 ;
        RECT 108.535 119.105 108.790 119.675 ;
        RECT 109.340 119.645 109.520 120.295 ;
        RECT 110.240 120.175 110.490 120.765 ;
        RECT 110.840 120.615 111.010 121.225 ;
        RECT 111.180 120.795 111.510 121.485 ;
        RECT 111.740 120.935 111.980 121.225 ;
        RECT 112.180 121.105 112.600 121.485 ;
        RECT 112.780 121.015 113.410 121.265 ;
        RECT 113.880 121.105 114.210 121.485 ;
        RECT 112.780 120.935 112.950 121.015 ;
        RECT 114.380 120.935 114.550 121.225 ;
        RECT 114.730 121.105 115.110 121.485 ;
        RECT 115.350 121.100 116.180 121.270 ;
        RECT 111.740 120.765 112.950 120.935 ;
        RECT 109.690 119.845 110.490 120.175 ;
        RECT 109.340 119.115 109.595 119.645 ;
        RECT 109.775 118.935 110.060 119.395 ;
        RECT 110.240 119.195 110.490 119.845 ;
        RECT 110.690 120.595 111.010 120.615 ;
        RECT 110.690 120.425 112.610 120.595 ;
        RECT 110.690 119.530 110.880 120.425 ;
        RECT 112.780 120.255 112.950 120.765 ;
        RECT 113.120 120.505 113.640 120.815 ;
        RECT 111.050 120.085 112.950 120.255 ;
        RECT 111.050 120.025 111.380 120.085 ;
        RECT 111.530 119.855 111.860 119.915 ;
        RECT 111.200 119.585 111.860 119.855 ;
        RECT 110.690 119.200 111.010 119.530 ;
        RECT 111.190 118.935 111.850 119.415 ;
        RECT 112.050 119.325 112.220 120.085 ;
        RECT 113.120 119.915 113.300 120.325 ;
        RECT 112.390 119.745 112.720 119.865 ;
        RECT 113.470 119.745 113.640 120.505 ;
        RECT 112.390 119.575 113.640 119.745 ;
        RECT 113.810 120.685 115.180 120.935 ;
        RECT 113.810 119.915 114.000 120.685 ;
        RECT 114.930 120.425 115.180 120.685 ;
        RECT 114.170 120.255 114.420 120.415 ;
        RECT 115.350 120.255 115.520 121.100 ;
        RECT 116.415 120.815 116.585 121.315 ;
        RECT 116.755 120.985 117.085 121.485 ;
        RECT 115.690 120.425 116.190 120.805 ;
        RECT 116.415 120.645 117.110 120.815 ;
        RECT 114.170 120.085 115.520 120.255 ;
        RECT 115.100 120.045 115.520 120.085 ;
        RECT 113.810 119.575 114.230 119.915 ;
        RECT 114.520 119.585 114.930 119.915 ;
        RECT 112.050 119.155 112.900 119.325 ;
        RECT 113.460 118.935 113.780 119.395 ;
        RECT 113.980 119.145 114.230 119.575 ;
        RECT 114.520 118.935 114.930 119.375 ;
        RECT 115.100 119.315 115.270 120.045 ;
        RECT 115.440 119.495 115.790 119.865 ;
        RECT 115.970 119.555 116.190 120.425 ;
        RECT 116.360 119.855 116.770 120.475 ;
        RECT 116.940 119.675 117.110 120.645 ;
        RECT 116.415 119.485 117.110 119.675 ;
        RECT 115.100 119.115 116.115 119.315 ;
        RECT 116.415 119.155 116.585 119.485 ;
        RECT 116.755 118.935 117.085 119.315 ;
        RECT 117.300 119.195 117.525 121.315 ;
        RECT 117.695 120.985 118.025 121.485 ;
        RECT 118.195 120.815 118.365 121.315 ;
        RECT 117.700 120.645 118.365 120.815 ;
        RECT 117.700 119.655 117.930 120.645 ;
        RECT 118.100 119.825 118.450 120.475 ;
        RECT 118.665 120.345 118.895 121.485 ;
        RECT 119.065 120.335 119.395 121.315 ;
        RECT 119.565 120.345 119.775 121.485 ;
        RECT 120.555 120.555 120.725 121.315 ;
        RECT 120.905 120.725 121.235 121.485 ;
        RECT 120.555 120.385 121.220 120.555 ;
        RECT 121.405 120.410 121.675 121.315 ;
        RECT 118.645 119.925 118.975 120.175 ;
        RECT 117.700 119.485 118.365 119.655 ;
        RECT 117.695 118.935 118.025 119.315 ;
        RECT 118.195 119.195 118.365 119.485 ;
        RECT 118.665 118.935 118.895 119.755 ;
        RECT 119.145 119.735 119.395 120.335 ;
        RECT 121.050 120.240 121.220 120.385 ;
        RECT 120.485 119.835 120.815 120.205 ;
        RECT 121.050 119.910 121.335 120.240 ;
        RECT 119.065 119.105 119.395 119.735 ;
        RECT 119.565 118.935 119.775 119.755 ;
        RECT 121.050 119.655 121.220 119.910 ;
        RECT 120.555 119.485 121.220 119.655 ;
        RECT 121.505 119.610 121.675 120.410 ;
        RECT 122.765 120.395 126.275 121.485 ;
        RECT 126.445 120.395 127.655 121.485 ;
        RECT 122.765 119.875 124.455 120.395 ;
        RECT 124.625 119.705 126.275 120.225 ;
        RECT 126.445 119.855 126.965 120.395 ;
        RECT 120.555 119.105 120.725 119.485 ;
        RECT 120.905 118.935 121.235 119.315 ;
        RECT 121.415 119.105 121.675 119.610 ;
        RECT 122.765 118.935 126.275 119.705 ;
        RECT 127.135 119.685 127.655 120.225 ;
        RECT 126.445 118.935 127.655 119.685 ;
        RECT 14.580 118.765 127.740 118.935 ;
        RECT 14.665 118.015 15.875 118.765 ;
        RECT 14.665 117.475 15.185 118.015 ;
        RECT 16.565 117.945 16.775 118.765 ;
        RECT 16.945 117.965 17.275 118.595 ;
        RECT 15.355 117.305 15.875 117.845 ;
        RECT 16.945 117.365 17.195 117.965 ;
        RECT 17.445 117.945 17.675 118.765 ;
        RECT 18.260 118.425 18.515 118.585 ;
        RECT 18.175 118.255 18.515 118.425 ;
        RECT 18.695 118.305 18.980 118.765 ;
        RECT 18.260 118.055 18.515 118.255 ;
        RECT 17.365 117.525 17.695 117.775 ;
        RECT 14.665 116.215 15.875 117.305 ;
        RECT 16.565 116.215 16.775 117.355 ;
        RECT 16.945 116.385 17.275 117.365 ;
        RECT 17.445 116.215 17.675 117.355 ;
        RECT 18.260 117.195 18.440 118.055 ;
        RECT 19.160 117.855 19.410 118.505 ;
        RECT 18.610 117.525 19.410 117.855 ;
        RECT 18.260 116.525 18.515 117.195 ;
        RECT 18.695 116.215 18.980 117.015 ;
        RECT 19.160 116.935 19.410 117.525 ;
        RECT 19.610 118.170 19.930 118.500 ;
        RECT 20.110 118.285 20.770 118.765 ;
        RECT 20.970 118.375 21.820 118.545 ;
        RECT 19.610 117.275 19.800 118.170 ;
        RECT 20.120 117.845 20.780 118.115 ;
        RECT 20.450 117.785 20.780 117.845 ;
        RECT 19.970 117.615 20.300 117.675 ;
        RECT 20.970 117.615 21.140 118.375 ;
        RECT 22.380 118.305 22.700 118.765 ;
        RECT 22.900 118.125 23.150 118.555 ;
        RECT 23.440 118.325 23.850 118.765 ;
        RECT 24.020 118.385 25.035 118.585 ;
        RECT 21.310 117.955 22.560 118.125 ;
        RECT 21.310 117.835 21.640 117.955 ;
        RECT 19.970 117.445 21.870 117.615 ;
        RECT 19.610 117.105 21.530 117.275 ;
        RECT 19.610 117.085 19.930 117.105 ;
        RECT 19.160 116.425 19.490 116.935 ;
        RECT 19.760 116.475 19.930 117.085 ;
        RECT 21.700 116.935 21.870 117.445 ;
        RECT 22.040 117.375 22.220 117.785 ;
        RECT 22.390 117.195 22.560 117.955 ;
        RECT 20.100 116.215 20.430 116.905 ;
        RECT 20.660 116.765 21.870 116.935 ;
        RECT 22.040 116.885 22.560 117.195 ;
        RECT 22.730 117.785 23.150 118.125 ;
        RECT 23.440 117.785 23.850 118.115 ;
        RECT 22.730 117.015 22.920 117.785 ;
        RECT 24.020 117.655 24.190 118.385 ;
        RECT 25.335 118.215 25.505 118.545 ;
        RECT 25.675 118.385 26.005 118.765 ;
        RECT 24.360 117.835 24.710 118.205 ;
        RECT 24.020 117.615 24.440 117.655 ;
        RECT 23.090 117.445 24.440 117.615 ;
        RECT 23.090 117.285 23.340 117.445 ;
        RECT 23.850 117.015 24.100 117.275 ;
        RECT 22.730 116.765 24.100 117.015 ;
        RECT 20.660 116.475 20.900 116.765 ;
        RECT 21.700 116.685 21.870 116.765 ;
        RECT 21.100 116.215 21.520 116.595 ;
        RECT 21.700 116.435 22.330 116.685 ;
        RECT 22.800 116.215 23.130 116.595 ;
        RECT 23.300 116.475 23.470 116.765 ;
        RECT 24.270 116.600 24.440 117.445 ;
        RECT 24.890 117.275 25.110 118.145 ;
        RECT 25.335 118.025 26.030 118.215 ;
        RECT 24.610 116.895 25.110 117.275 ;
        RECT 25.280 117.225 25.690 117.845 ;
        RECT 25.860 117.055 26.030 118.025 ;
        RECT 25.335 116.885 26.030 117.055 ;
        RECT 23.650 116.215 24.030 116.595 ;
        RECT 24.270 116.430 25.100 116.600 ;
        RECT 25.335 116.385 25.505 116.885 ;
        RECT 25.675 116.215 26.005 116.715 ;
        RECT 26.220 116.385 26.445 118.505 ;
        RECT 26.615 118.385 26.945 118.765 ;
        RECT 27.115 118.215 27.285 118.505 ;
        RECT 26.620 118.045 27.285 118.215 ;
        RECT 27.635 118.215 27.805 118.505 ;
        RECT 27.975 118.385 28.305 118.765 ;
        RECT 27.635 118.045 28.300 118.215 ;
        RECT 26.620 117.055 26.850 118.045 ;
        RECT 27.020 117.225 27.370 117.875 ;
        RECT 27.550 117.225 27.900 117.875 ;
        RECT 28.070 117.055 28.300 118.045 ;
        RECT 26.620 116.885 27.285 117.055 ;
        RECT 26.615 116.215 26.945 116.715 ;
        RECT 27.115 116.385 27.285 116.885 ;
        RECT 27.635 116.885 28.300 117.055 ;
        RECT 27.635 116.385 27.805 116.885 ;
        RECT 27.975 116.215 28.305 116.715 ;
        RECT 28.475 116.385 28.700 118.505 ;
        RECT 28.915 118.385 29.245 118.765 ;
        RECT 29.415 118.215 29.585 118.545 ;
        RECT 29.885 118.385 30.900 118.585 ;
        RECT 28.890 118.025 29.585 118.215 ;
        RECT 28.890 117.055 29.060 118.025 ;
        RECT 29.230 117.225 29.640 117.845 ;
        RECT 29.810 117.275 30.030 118.145 ;
        RECT 30.210 117.835 30.560 118.205 ;
        RECT 30.730 117.655 30.900 118.385 ;
        RECT 31.070 118.325 31.480 118.765 ;
        RECT 31.770 118.125 32.020 118.555 ;
        RECT 32.220 118.305 32.540 118.765 ;
        RECT 33.100 118.375 33.950 118.545 ;
        RECT 31.070 117.785 31.480 118.115 ;
        RECT 31.770 117.785 32.190 118.125 ;
        RECT 30.480 117.615 30.900 117.655 ;
        RECT 30.480 117.445 31.830 117.615 ;
        RECT 28.890 116.885 29.585 117.055 ;
        RECT 29.810 116.895 30.310 117.275 ;
        RECT 28.915 116.215 29.245 116.715 ;
        RECT 29.415 116.385 29.585 116.885 ;
        RECT 30.480 116.600 30.650 117.445 ;
        RECT 31.580 117.285 31.830 117.445 ;
        RECT 30.820 117.015 31.070 117.275 ;
        RECT 32.000 117.015 32.190 117.785 ;
        RECT 30.820 116.765 32.190 117.015 ;
        RECT 32.360 117.955 33.610 118.125 ;
        RECT 32.360 117.195 32.530 117.955 ;
        RECT 33.280 117.835 33.610 117.955 ;
        RECT 32.700 117.375 32.880 117.785 ;
        RECT 33.780 117.615 33.950 118.375 ;
        RECT 34.150 118.285 34.810 118.765 ;
        RECT 34.990 118.170 35.310 118.500 ;
        RECT 34.140 117.845 34.800 118.115 ;
        RECT 34.140 117.785 34.470 117.845 ;
        RECT 34.620 117.615 34.950 117.675 ;
        RECT 33.050 117.445 34.950 117.615 ;
        RECT 32.360 116.885 32.880 117.195 ;
        RECT 33.050 116.935 33.220 117.445 ;
        RECT 35.120 117.275 35.310 118.170 ;
        RECT 33.390 117.105 35.310 117.275 ;
        RECT 34.990 117.085 35.310 117.105 ;
        RECT 35.510 117.855 35.760 118.505 ;
        RECT 35.940 118.305 36.225 118.765 ;
        RECT 36.405 118.425 36.660 118.585 ;
        RECT 36.405 118.255 36.745 118.425 ;
        RECT 36.405 118.055 36.660 118.255 ;
        RECT 35.510 117.525 36.310 117.855 ;
        RECT 33.050 116.765 34.260 116.935 ;
        RECT 29.820 116.430 30.650 116.600 ;
        RECT 30.890 116.215 31.270 116.595 ;
        RECT 31.450 116.475 31.620 116.765 ;
        RECT 33.050 116.685 33.220 116.765 ;
        RECT 31.790 116.215 32.120 116.595 ;
        RECT 32.590 116.435 33.220 116.685 ;
        RECT 33.400 116.215 33.820 116.595 ;
        RECT 34.020 116.475 34.260 116.765 ;
        RECT 34.490 116.215 34.820 116.905 ;
        RECT 34.990 116.475 35.160 117.085 ;
        RECT 35.510 116.935 35.760 117.525 ;
        RECT 36.480 117.195 36.660 118.055 ;
        RECT 37.205 118.040 37.495 118.765 ;
        RECT 38.040 118.425 38.295 118.585 ;
        RECT 37.955 118.255 38.295 118.425 ;
        RECT 38.475 118.305 38.760 118.765 ;
        RECT 38.040 118.055 38.295 118.255 ;
        RECT 35.430 116.425 35.760 116.935 ;
        RECT 35.940 116.215 36.225 117.015 ;
        RECT 36.405 116.525 36.660 117.195 ;
        RECT 37.205 116.215 37.495 117.380 ;
        RECT 38.040 117.195 38.220 118.055 ;
        RECT 38.940 117.855 39.190 118.505 ;
        RECT 38.390 117.525 39.190 117.855 ;
        RECT 38.040 116.525 38.295 117.195 ;
        RECT 38.475 116.215 38.760 117.015 ;
        RECT 38.940 116.935 39.190 117.525 ;
        RECT 39.390 118.170 39.710 118.500 ;
        RECT 39.890 118.285 40.550 118.765 ;
        RECT 40.750 118.375 41.600 118.545 ;
        RECT 39.390 117.275 39.580 118.170 ;
        RECT 39.900 117.845 40.560 118.115 ;
        RECT 40.230 117.785 40.560 117.845 ;
        RECT 39.750 117.615 40.080 117.675 ;
        RECT 40.750 117.615 40.920 118.375 ;
        RECT 42.160 118.305 42.480 118.765 ;
        RECT 42.680 118.125 42.930 118.555 ;
        RECT 43.220 118.325 43.630 118.765 ;
        RECT 43.800 118.385 44.815 118.585 ;
        RECT 41.090 117.955 42.340 118.125 ;
        RECT 41.090 117.835 41.420 117.955 ;
        RECT 39.750 117.445 41.650 117.615 ;
        RECT 39.390 117.105 41.310 117.275 ;
        RECT 39.390 117.085 39.710 117.105 ;
        RECT 38.940 116.425 39.270 116.935 ;
        RECT 39.540 116.475 39.710 117.085 ;
        RECT 41.480 116.935 41.650 117.445 ;
        RECT 41.820 117.375 42.000 117.785 ;
        RECT 42.170 117.195 42.340 117.955 ;
        RECT 39.880 116.215 40.210 116.905 ;
        RECT 40.440 116.765 41.650 116.935 ;
        RECT 41.820 116.885 42.340 117.195 ;
        RECT 42.510 117.785 42.930 118.125 ;
        RECT 43.220 117.785 43.630 118.115 ;
        RECT 42.510 117.015 42.700 117.785 ;
        RECT 43.800 117.655 43.970 118.385 ;
        RECT 45.115 118.215 45.285 118.545 ;
        RECT 45.455 118.385 45.785 118.765 ;
        RECT 44.140 117.835 44.490 118.205 ;
        RECT 43.800 117.615 44.220 117.655 ;
        RECT 42.870 117.445 44.220 117.615 ;
        RECT 42.870 117.285 43.120 117.445 ;
        RECT 43.630 117.015 43.880 117.275 ;
        RECT 42.510 116.765 43.880 117.015 ;
        RECT 40.440 116.475 40.680 116.765 ;
        RECT 41.480 116.685 41.650 116.765 ;
        RECT 40.880 116.215 41.300 116.595 ;
        RECT 41.480 116.435 42.110 116.685 ;
        RECT 42.580 116.215 42.910 116.595 ;
        RECT 43.080 116.475 43.250 116.765 ;
        RECT 44.050 116.600 44.220 117.445 ;
        RECT 44.670 117.275 44.890 118.145 ;
        RECT 45.115 118.025 45.810 118.215 ;
        RECT 44.390 116.895 44.890 117.275 ;
        RECT 45.060 117.225 45.470 117.845 ;
        RECT 45.640 117.055 45.810 118.025 ;
        RECT 45.115 116.885 45.810 117.055 ;
        RECT 43.430 116.215 43.810 116.595 ;
        RECT 44.050 116.430 44.880 116.600 ;
        RECT 45.115 116.385 45.285 116.885 ;
        RECT 45.455 116.215 45.785 116.715 ;
        RECT 46.000 116.385 46.225 118.505 ;
        RECT 46.395 118.385 46.725 118.765 ;
        RECT 46.895 118.215 47.065 118.505 ;
        RECT 46.400 118.045 47.065 118.215 ;
        RECT 47.700 118.055 47.955 118.585 ;
        RECT 48.135 118.305 48.420 118.765 ;
        RECT 46.400 117.055 46.630 118.045 ;
        RECT 46.800 117.225 47.150 117.875 ;
        RECT 47.700 117.195 47.880 118.055 ;
        RECT 48.600 117.855 48.850 118.505 ;
        RECT 48.050 117.525 48.850 117.855 ;
        RECT 46.400 116.885 47.065 117.055 ;
        RECT 46.395 116.215 46.725 116.715 ;
        RECT 46.895 116.385 47.065 116.885 ;
        RECT 47.700 116.725 47.955 117.195 ;
        RECT 47.615 116.555 47.955 116.725 ;
        RECT 47.700 116.525 47.955 116.555 ;
        RECT 48.135 116.215 48.420 117.015 ;
        RECT 48.600 116.935 48.850 117.525 ;
        RECT 49.050 118.170 49.370 118.500 ;
        RECT 49.550 118.285 50.210 118.765 ;
        RECT 50.410 118.375 51.260 118.545 ;
        RECT 49.050 117.275 49.240 118.170 ;
        RECT 49.560 117.845 50.220 118.115 ;
        RECT 49.890 117.785 50.220 117.845 ;
        RECT 49.410 117.615 49.740 117.675 ;
        RECT 50.410 117.615 50.580 118.375 ;
        RECT 51.820 118.305 52.140 118.765 ;
        RECT 52.340 118.125 52.590 118.555 ;
        RECT 52.880 118.325 53.290 118.765 ;
        RECT 53.460 118.385 54.475 118.585 ;
        RECT 50.750 117.955 52.000 118.125 ;
        RECT 50.750 117.835 51.080 117.955 ;
        RECT 49.410 117.445 51.310 117.615 ;
        RECT 49.050 117.105 50.970 117.275 ;
        RECT 49.050 117.085 49.370 117.105 ;
        RECT 48.600 116.425 48.930 116.935 ;
        RECT 49.200 116.475 49.370 117.085 ;
        RECT 51.140 116.935 51.310 117.445 ;
        RECT 51.480 117.375 51.660 117.785 ;
        RECT 51.830 117.195 52.000 117.955 ;
        RECT 49.540 116.215 49.870 116.905 ;
        RECT 50.100 116.765 51.310 116.935 ;
        RECT 51.480 116.885 52.000 117.195 ;
        RECT 52.170 117.785 52.590 118.125 ;
        RECT 52.880 117.785 53.290 118.115 ;
        RECT 52.170 117.015 52.360 117.785 ;
        RECT 53.460 117.655 53.630 118.385 ;
        RECT 54.775 118.215 54.945 118.545 ;
        RECT 55.115 118.385 55.445 118.765 ;
        RECT 53.800 117.835 54.150 118.205 ;
        RECT 53.460 117.615 53.880 117.655 ;
        RECT 52.530 117.445 53.880 117.615 ;
        RECT 52.530 117.285 52.780 117.445 ;
        RECT 53.290 117.015 53.540 117.275 ;
        RECT 52.170 116.765 53.540 117.015 ;
        RECT 50.100 116.475 50.340 116.765 ;
        RECT 51.140 116.685 51.310 116.765 ;
        RECT 50.540 116.215 50.960 116.595 ;
        RECT 51.140 116.435 51.770 116.685 ;
        RECT 52.240 116.215 52.570 116.595 ;
        RECT 52.740 116.475 52.910 116.765 ;
        RECT 53.710 116.600 53.880 117.445 ;
        RECT 54.330 117.275 54.550 118.145 ;
        RECT 54.775 118.025 55.470 118.215 ;
        RECT 54.050 116.895 54.550 117.275 ;
        RECT 54.720 117.225 55.130 117.845 ;
        RECT 55.300 117.055 55.470 118.025 ;
        RECT 54.775 116.885 55.470 117.055 ;
        RECT 53.090 116.215 53.470 116.595 ;
        RECT 53.710 116.430 54.540 116.600 ;
        RECT 54.775 116.385 54.945 116.885 ;
        RECT 55.115 116.215 55.445 116.715 ;
        RECT 55.660 116.385 55.885 118.505 ;
        RECT 56.055 118.385 56.385 118.765 ;
        RECT 56.555 118.215 56.725 118.505 ;
        RECT 56.060 118.045 56.725 118.215 ;
        RECT 56.060 117.055 56.290 118.045 ;
        RECT 57.905 117.995 61.415 118.765 ;
        RECT 56.460 117.225 56.810 117.875 ;
        RECT 57.905 117.305 59.595 117.825 ;
        RECT 59.765 117.475 61.415 117.995 ;
        RECT 61.625 117.945 61.855 118.765 ;
        RECT 62.025 117.965 62.355 118.595 ;
        RECT 61.605 117.525 61.935 117.775 ;
        RECT 62.105 117.365 62.355 117.965 ;
        RECT 62.525 117.945 62.735 118.765 ;
        RECT 62.965 118.040 63.255 118.765 ;
        RECT 63.800 118.425 64.055 118.585 ;
        RECT 63.715 118.255 64.055 118.425 ;
        RECT 64.235 118.305 64.520 118.765 ;
        RECT 63.800 118.055 64.055 118.255 ;
        RECT 56.060 116.885 56.725 117.055 ;
        RECT 56.055 116.215 56.385 116.715 ;
        RECT 56.555 116.385 56.725 116.885 ;
        RECT 57.905 116.215 61.415 117.305 ;
        RECT 61.625 116.215 61.855 117.355 ;
        RECT 62.025 116.385 62.355 117.365 ;
        RECT 62.525 116.215 62.735 117.355 ;
        RECT 62.965 116.215 63.255 117.380 ;
        RECT 63.800 117.195 63.980 118.055 ;
        RECT 64.700 117.855 64.950 118.505 ;
        RECT 64.150 117.525 64.950 117.855 ;
        RECT 63.800 116.525 64.055 117.195 ;
        RECT 64.235 116.215 64.520 117.015 ;
        RECT 64.700 116.935 64.950 117.525 ;
        RECT 65.150 118.170 65.470 118.500 ;
        RECT 65.650 118.285 66.310 118.765 ;
        RECT 66.510 118.375 67.360 118.545 ;
        RECT 65.150 117.275 65.340 118.170 ;
        RECT 65.660 117.845 66.320 118.115 ;
        RECT 65.990 117.785 66.320 117.845 ;
        RECT 65.510 117.615 65.840 117.675 ;
        RECT 66.510 117.615 66.680 118.375 ;
        RECT 67.920 118.305 68.240 118.765 ;
        RECT 68.440 118.125 68.690 118.555 ;
        RECT 68.980 118.325 69.390 118.765 ;
        RECT 69.560 118.385 70.575 118.585 ;
        RECT 66.850 117.955 68.100 118.125 ;
        RECT 66.850 117.835 67.180 117.955 ;
        RECT 65.510 117.445 67.410 117.615 ;
        RECT 65.150 117.105 67.070 117.275 ;
        RECT 65.150 117.085 65.470 117.105 ;
        RECT 64.700 116.425 65.030 116.935 ;
        RECT 65.300 116.475 65.470 117.085 ;
        RECT 67.240 116.935 67.410 117.445 ;
        RECT 67.580 117.375 67.760 117.785 ;
        RECT 67.930 117.195 68.100 117.955 ;
        RECT 65.640 116.215 65.970 116.905 ;
        RECT 66.200 116.765 67.410 116.935 ;
        RECT 67.580 116.885 68.100 117.195 ;
        RECT 68.270 117.785 68.690 118.125 ;
        RECT 68.980 117.785 69.390 118.115 ;
        RECT 68.270 117.015 68.460 117.785 ;
        RECT 69.560 117.655 69.730 118.385 ;
        RECT 70.875 118.215 71.045 118.545 ;
        RECT 71.215 118.385 71.545 118.765 ;
        RECT 69.900 117.835 70.250 118.205 ;
        RECT 69.560 117.615 69.980 117.655 ;
        RECT 68.630 117.445 69.980 117.615 ;
        RECT 68.630 117.285 68.880 117.445 ;
        RECT 69.390 117.015 69.640 117.275 ;
        RECT 68.270 116.765 69.640 117.015 ;
        RECT 66.200 116.475 66.440 116.765 ;
        RECT 67.240 116.685 67.410 116.765 ;
        RECT 66.640 116.215 67.060 116.595 ;
        RECT 67.240 116.435 67.870 116.685 ;
        RECT 68.340 116.215 68.670 116.595 ;
        RECT 68.840 116.475 69.010 116.765 ;
        RECT 69.810 116.600 69.980 117.445 ;
        RECT 70.430 117.275 70.650 118.145 ;
        RECT 70.875 118.025 71.570 118.215 ;
        RECT 70.150 116.895 70.650 117.275 ;
        RECT 70.820 117.225 71.230 117.845 ;
        RECT 71.400 117.055 71.570 118.025 ;
        RECT 70.875 116.885 71.570 117.055 ;
        RECT 69.190 116.215 69.570 116.595 ;
        RECT 69.810 116.430 70.640 116.600 ;
        RECT 70.875 116.385 71.045 116.885 ;
        RECT 71.215 116.215 71.545 116.715 ;
        RECT 71.760 116.385 71.985 118.505 ;
        RECT 72.155 118.385 72.485 118.765 ;
        RECT 72.655 118.215 72.825 118.505 ;
        RECT 73.460 118.425 73.715 118.585 ;
        RECT 73.375 118.255 73.715 118.425 ;
        RECT 73.895 118.305 74.180 118.765 ;
        RECT 72.160 118.045 72.825 118.215 ;
        RECT 73.460 118.055 73.715 118.255 ;
        RECT 72.160 117.055 72.390 118.045 ;
        RECT 72.560 117.225 72.910 117.875 ;
        RECT 73.460 117.195 73.640 118.055 ;
        RECT 74.360 117.855 74.610 118.505 ;
        RECT 73.810 117.525 74.610 117.855 ;
        RECT 72.160 116.885 72.825 117.055 ;
        RECT 72.155 116.215 72.485 116.715 ;
        RECT 72.655 116.385 72.825 116.885 ;
        RECT 73.460 116.525 73.715 117.195 ;
        RECT 73.895 116.215 74.180 117.015 ;
        RECT 74.360 116.935 74.610 117.525 ;
        RECT 74.810 118.170 75.130 118.500 ;
        RECT 75.310 118.285 75.970 118.765 ;
        RECT 76.170 118.375 77.020 118.545 ;
        RECT 74.810 117.275 75.000 118.170 ;
        RECT 75.320 117.845 75.980 118.115 ;
        RECT 75.650 117.785 75.980 117.845 ;
        RECT 75.170 117.615 75.500 117.675 ;
        RECT 76.170 117.615 76.340 118.375 ;
        RECT 77.580 118.305 77.900 118.765 ;
        RECT 78.100 118.125 78.350 118.555 ;
        RECT 78.640 118.325 79.050 118.765 ;
        RECT 79.220 118.385 80.235 118.585 ;
        RECT 76.510 117.955 77.760 118.125 ;
        RECT 76.510 117.835 76.840 117.955 ;
        RECT 75.170 117.445 77.070 117.615 ;
        RECT 74.810 117.105 76.730 117.275 ;
        RECT 74.810 117.085 75.130 117.105 ;
        RECT 74.360 116.425 74.690 116.935 ;
        RECT 74.960 116.475 75.130 117.085 ;
        RECT 76.900 116.935 77.070 117.445 ;
        RECT 77.240 117.375 77.420 117.785 ;
        RECT 77.590 117.195 77.760 117.955 ;
        RECT 75.300 116.215 75.630 116.905 ;
        RECT 75.860 116.765 77.070 116.935 ;
        RECT 77.240 116.885 77.760 117.195 ;
        RECT 77.930 117.785 78.350 118.125 ;
        RECT 78.640 117.785 79.050 118.115 ;
        RECT 77.930 117.015 78.120 117.785 ;
        RECT 79.220 117.655 79.390 118.385 ;
        RECT 80.535 118.215 80.705 118.545 ;
        RECT 80.875 118.385 81.205 118.765 ;
        RECT 79.560 117.835 79.910 118.205 ;
        RECT 79.220 117.615 79.640 117.655 ;
        RECT 78.290 117.445 79.640 117.615 ;
        RECT 78.290 117.285 78.540 117.445 ;
        RECT 79.050 117.015 79.300 117.275 ;
        RECT 77.930 116.765 79.300 117.015 ;
        RECT 75.860 116.475 76.100 116.765 ;
        RECT 76.900 116.685 77.070 116.765 ;
        RECT 76.300 116.215 76.720 116.595 ;
        RECT 76.900 116.435 77.530 116.685 ;
        RECT 78.000 116.215 78.330 116.595 ;
        RECT 78.500 116.475 78.670 116.765 ;
        RECT 79.470 116.600 79.640 117.445 ;
        RECT 80.090 117.275 80.310 118.145 ;
        RECT 80.535 118.025 81.230 118.215 ;
        RECT 79.810 116.895 80.310 117.275 ;
        RECT 80.480 117.225 80.890 117.845 ;
        RECT 81.060 117.055 81.230 118.025 ;
        RECT 80.535 116.885 81.230 117.055 ;
        RECT 78.850 116.215 79.230 116.595 ;
        RECT 79.470 116.430 80.300 116.600 ;
        RECT 80.535 116.385 80.705 116.885 ;
        RECT 80.875 116.215 81.205 116.715 ;
        RECT 81.420 116.385 81.645 118.505 ;
        RECT 81.815 118.385 82.145 118.765 ;
        RECT 82.315 118.215 82.485 118.505 ;
        RECT 81.820 118.045 82.485 118.215 ;
        RECT 81.820 117.055 82.050 118.045 ;
        RECT 82.750 118.025 83.005 118.595 ;
        RECT 83.175 118.365 83.505 118.765 ;
        RECT 83.930 118.230 84.460 118.595 ;
        RECT 83.930 118.195 84.105 118.230 ;
        RECT 83.175 118.025 84.105 118.195 ;
        RECT 82.220 117.225 82.570 117.875 ;
        RECT 82.750 117.355 82.920 118.025 ;
        RECT 83.175 117.855 83.345 118.025 ;
        RECT 83.090 117.525 83.345 117.855 ;
        RECT 83.570 117.525 83.765 117.855 ;
        RECT 81.820 116.885 82.485 117.055 ;
        RECT 81.815 116.215 82.145 116.715 ;
        RECT 82.315 116.385 82.485 116.885 ;
        RECT 82.750 116.385 83.085 117.355 ;
        RECT 83.255 116.215 83.425 117.355 ;
        RECT 83.595 116.555 83.765 117.525 ;
        RECT 83.935 116.895 84.105 118.025 ;
        RECT 84.275 117.235 84.445 118.035 ;
        RECT 84.650 117.745 84.925 118.595 ;
        RECT 84.645 117.575 84.925 117.745 ;
        RECT 84.650 117.435 84.925 117.575 ;
        RECT 85.095 117.235 85.285 118.595 ;
        RECT 85.465 118.230 85.975 118.765 ;
        RECT 86.195 117.955 86.440 118.560 ;
        RECT 87.435 118.215 87.605 118.595 ;
        RECT 87.785 118.385 88.115 118.765 ;
        RECT 87.435 118.045 88.100 118.215 ;
        RECT 88.295 118.090 88.555 118.595 ;
        RECT 85.485 117.785 86.715 117.955 ;
        RECT 84.275 117.065 85.285 117.235 ;
        RECT 85.455 117.220 86.205 117.410 ;
        RECT 83.935 116.725 85.060 116.895 ;
        RECT 85.455 116.555 85.625 117.220 ;
        RECT 86.375 116.975 86.715 117.785 ;
        RECT 87.365 117.495 87.695 117.865 ;
        RECT 87.930 117.790 88.100 118.045 ;
        RECT 87.930 117.460 88.215 117.790 ;
        RECT 87.930 117.315 88.100 117.460 ;
        RECT 83.595 116.385 85.625 116.555 ;
        RECT 85.795 116.215 85.965 116.975 ;
        RECT 86.200 116.565 86.715 116.975 ;
        RECT 87.435 117.145 88.100 117.315 ;
        RECT 88.385 117.290 88.555 118.090 ;
        RECT 88.725 118.040 89.015 118.765 ;
        RECT 89.225 117.945 89.455 118.765 ;
        RECT 89.625 117.965 89.955 118.595 ;
        RECT 89.205 117.525 89.535 117.775 ;
        RECT 87.435 116.385 87.605 117.145 ;
        RECT 87.785 116.215 88.115 116.975 ;
        RECT 88.285 116.385 88.555 117.290 ;
        RECT 88.725 116.215 89.015 117.380 ;
        RECT 89.705 117.365 89.955 117.965 ;
        RECT 90.125 117.945 90.335 118.765 ;
        RECT 90.605 117.945 90.835 118.765 ;
        RECT 91.005 117.965 91.335 118.595 ;
        RECT 90.585 117.525 90.915 117.775 ;
        RECT 91.085 117.365 91.335 117.965 ;
        RECT 91.505 117.945 91.715 118.765 ;
        RECT 93.240 118.425 93.495 118.585 ;
        RECT 93.155 118.255 93.495 118.425 ;
        RECT 93.675 118.305 93.960 118.765 ;
        RECT 93.240 118.055 93.495 118.255 ;
        RECT 89.225 116.215 89.455 117.355 ;
        RECT 89.625 116.385 89.955 117.365 ;
        RECT 90.125 116.215 90.335 117.355 ;
        RECT 90.605 116.215 90.835 117.355 ;
        RECT 91.005 116.385 91.335 117.365 ;
        RECT 91.505 116.215 91.715 117.355 ;
        RECT 93.240 117.195 93.420 118.055 ;
        RECT 94.140 117.855 94.390 118.505 ;
        RECT 93.590 117.525 94.390 117.855 ;
        RECT 93.240 116.525 93.495 117.195 ;
        RECT 93.675 116.215 93.960 117.015 ;
        RECT 94.140 116.935 94.390 117.525 ;
        RECT 94.590 118.170 94.910 118.500 ;
        RECT 95.090 118.285 95.750 118.765 ;
        RECT 95.950 118.375 96.800 118.545 ;
        RECT 94.590 117.275 94.780 118.170 ;
        RECT 95.100 117.845 95.760 118.115 ;
        RECT 95.430 117.785 95.760 117.845 ;
        RECT 94.950 117.615 95.280 117.675 ;
        RECT 95.950 117.615 96.120 118.375 ;
        RECT 97.360 118.305 97.680 118.765 ;
        RECT 97.880 118.125 98.130 118.555 ;
        RECT 98.420 118.325 98.830 118.765 ;
        RECT 99.000 118.385 100.015 118.585 ;
        RECT 96.290 117.955 97.540 118.125 ;
        RECT 96.290 117.835 96.620 117.955 ;
        RECT 94.950 117.445 96.850 117.615 ;
        RECT 94.590 117.105 96.510 117.275 ;
        RECT 94.590 117.085 94.910 117.105 ;
        RECT 94.140 116.425 94.470 116.935 ;
        RECT 94.740 116.475 94.910 117.085 ;
        RECT 96.680 116.935 96.850 117.445 ;
        RECT 97.020 117.375 97.200 117.785 ;
        RECT 97.370 117.195 97.540 117.955 ;
        RECT 95.080 116.215 95.410 116.905 ;
        RECT 95.640 116.765 96.850 116.935 ;
        RECT 97.020 116.885 97.540 117.195 ;
        RECT 97.710 117.785 98.130 118.125 ;
        RECT 98.420 117.785 98.830 118.115 ;
        RECT 97.710 117.015 97.900 117.785 ;
        RECT 99.000 117.655 99.170 118.385 ;
        RECT 100.315 118.215 100.485 118.545 ;
        RECT 100.655 118.385 100.985 118.765 ;
        RECT 99.340 117.835 99.690 118.205 ;
        RECT 99.000 117.615 99.420 117.655 ;
        RECT 98.070 117.445 99.420 117.615 ;
        RECT 98.070 117.285 98.320 117.445 ;
        RECT 98.830 117.015 99.080 117.275 ;
        RECT 97.710 116.765 99.080 117.015 ;
        RECT 95.640 116.475 95.880 116.765 ;
        RECT 96.680 116.685 96.850 116.765 ;
        RECT 96.080 116.215 96.500 116.595 ;
        RECT 96.680 116.435 97.310 116.685 ;
        RECT 97.780 116.215 98.110 116.595 ;
        RECT 98.280 116.475 98.450 116.765 ;
        RECT 99.250 116.600 99.420 117.445 ;
        RECT 99.870 117.275 100.090 118.145 ;
        RECT 100.315 118.025 101.010 118.215 ;
        RECT 99.590 116.895 100.090 117.275 ;
        RECT 100.260 117.225 100.670 117.845 ;
        RECT 100.840 117.055 101.010 118.025 ;
        RECT 100.315 116.885 101.010 117.055 ;
        RECT 98.630 116.215 99.010 116.595 ;
        RECT 99.250 116.430 100.080 116.600 ;
        RECT 100.315 116.385 100.485 116.885 ;
        RECT 100.655 116.215 100.985 116.715 ;
        RECT 101.200 116.385 101.425 118.505 ;
        RECT 101.595 118.385 101.925 118.765 ;
        RECT 102.095 118.215 102.265 118.505 ;
        RECT 102.900 118.425 103.155 118.585 ;
        RECT 102.815 118.255 103.155 118.425 ;
        RECT 103.335 118.305 103.620 118.765 ;
        RECT 101.600 118.045 102.265 118.215 ;
        RECT 102.900 118.055 103.155 118.255 ;
        RECT 101.600 117.055 101.830 118.045 ;
        RECT 102.000 117.225 102.350 117.875 ;
        RECT 102.900 117.195 103.080 118.055 ;
        RECT 103.800 117.855 104.050 118.505 ;
        RECT 103.250 117.525 104.050 117.855 ;
        RECT 101.600 116.885 102.265 117.055 ;
        RECT 101.595 116.215 101.925 116.715 ;
        RECT 102.095 116.385 102.265 116.885 ;
        RECT 102.900 116.525 103.155 117.195 ;
        RECT 103.335 116.215 103.620 117.015 ;
        RECT 103.800 116.935 104.050 117.525 ;
        RECT 104.250 118.170 104.570 118.500 ;
        RECT 104.750 118.285 105.410 118.765 ;
        RECT 105.610 118.375 106.460 118.545 ;
        RECT 104.250 117.275 104.440 118.170 ;
        RECT 104.760 117.845 105.420 118.115 ;
        RECT 105.090 117.785 105.420 117.845 ;
        RECT 104.610 117.615 104.940 117.675 ;
        RECT 105.610 117.615 105.780 118.375 ;
        RECT 107.020 118.305 107.340 118.765 ;
        RECT 107.540 118.125 107.790 118.555 ;
        RECT 108.080 118.325 108.490 118.765 ;
        RECT 108.660 118.385 109.675 118.585 ;
        RECT 105.950 117.955 107.200 118.125 ;
        RECT 105.950 117.835 106.280 117.955 ;
        RECT 104.610 117.445 106.510 117.615 ;
        RECT 104.250 117.105 106.170 117.275 ;
        RECT 104.250 117.085 104.570 117.105 ;
        RECT 103.800 116.425 104.130 116.935 ;
        RECT 104.400 116.475 104.570 117.085 ;
        RECT 106.340 116.935 106.510 117.445 ;
        RECT 106.680 117.375 106.860 117.785 ;
        RECT 107.030 117.195 107.200 117.955 ;
        RECT 104.740 116.215 105.070 116.905 ;
        RECT 105.300 116.765 106.510 116.935 ;
        RECT 106.680 116.885 107.200 117.195 ;
        RECT 107.370 117.785 107.790 118.125 ;
        RECT 108.080 117.785 108.490 118.115 ;
        RECT 107.370 117.015 107.560 117.785 ;
        RECT 108.660 117.655 108.830 118.385 ;
        RECT 109.975 118.215 110.145 118.545 ;
        RECT 110.315 118.385 110.645 118.765 ;
        RECT 109.000 117.835 109.350 118.205 ;
        RECT 108.660 117.615 109.080 117.655 ;
        RECT 107.730 117.445 109.080 117.615 ;
        RECT 107.730 117.285 107.980 117.445 ;
        RECT 108.490 117.015 108.740 117.275 ;
        RECT 107.370 116.765 108.740 117.015 ;
        RECT 105.300 116.475 105.540 116.765 ;
        RECT 106.340 116.685 106.510 116.765 ;
        RECT 105.740 116.215 106.160 116.595 ;
        RECT 106.340 116.435 106.970 116.685 ;
        RECT 107.440 116.215 107.770 116.595 ;
        RECT 107.940 116.475 108.110 116.765 ;
        RECT 108.910 116.600 109.080 117.445 ;
        RECT 109.530 117.275 109.750 118.145 ;
        RECT 109.975 118.025 110.670 118.215 ;
        RECT 109.250 116.895 109.750 117.275 ;
        RECT 109.920 117.225 110.330 117.845 ;
        RECT 110.500 117.055 110.670 118.025 ;
        RECT 109.975 116.885 110.670 117.055 ;
        RECT 108.290 116.215 108.670 116.595 ;
        RECT 108.910 116.430 109.740 116.600 ;
        RECT 109.975 116.385 110.145 116.885 ;
        RECT 110.315 116.215 110.645 116.715 ;
        RECT 110.860 116.385 111.085 118.505 ;
        RECT 111.255 118.385 111.585 118.765 ;
        RECT 111.755 118.215 111.925 118.505 ;
        RECT 111.260 118.045 111.925 118.215 ;
        RECT 111.260 117.055 111.490 118.045 ;
        RECT 113.165 117.945 113.375 118.765 ;
        RECT 113.545 117.965 113.875 118.595 ;
        RECT 111.660 117.225 112.010 117.875 ;
        RECT 113.545 117.365 113.795 117.965 ;
        RECT 114.045 117.945 114.275 118.765 ;
        RECT 114.485 118.040 114.775 118.765 ;
        RECT 115.495 118.215 115.665 118.595 ;
        RECT 115.845 118.385 116.175 118.765 ;
        RECT 115.495 118.045 116.160 118.215 ;
        RECT 116.355 118.090 116.615 118.595 ;
        RECT 113.965 117.525 114.295 117.775 ;
        RECT 115.425 117.495 115.755 117.865 ;
        RECT 115.990 117.790 116.160 118.045 ;
        RECT 115.990 117.460 116.275 117.790 ;
        RECT 111.260 116.885 111.925 117.055 ;
        RECT 111.255 116.215 111.585 116.715 ;
        RECT 111.755 116.385 111.925 116.885 ;
        RECT 113.165 116.215 113.375 117.355 ;
        RECT 113.545 116.385 113.875 117.365 ;
        RECT 114.045 116.215 114.275 117.355 ;
        RECT 114.485 116.215 114.775 117.380 ;
        RECT 115.990 117.315 116.160 117.460 ;
        RECT 115.495 117.145 116.160 117.315 ;
        RECT 116.445 117.290 116.615 118.090 ;
        RECT 117.245 117.995 120.755 118.765 ;
        RECT 120.930 118.220 126.275 118.765 ;
        RECT 115.495 116.385 115.665 117.145 ;
        RECT 115.845 116.215 116.175 116.975 ;
        RECT 116.345 116.385 116.615 117.290 ;
        RECT 117.245 117.305 118.935 117.825 ;
        RECT 119.105 117.475 120.755 117.995 ;
        RECT 117.245 116.215 120.755 117.305 ;
        RECT 122.520 116.650 122.870 117.900 ;
        RECT 124.350 117.390 124.690 118.220 ;
        RECT 126.445 118.015 127.655 118.765 ;
        RECT 126.445 117.305 126.965 117.845 ;
        RECT 127.135 117.475 127.655 118.015 ;
        RECT 120.930 116.215 126.275 116.650 ;
        RECT 126.445 116.215 127.655 117.305 ;
        RECT 14.580 116.045 127.740 116.215 ;
        RECT 14.665 114.955 15.875 116.045 ;
        RECT 14.665 114.245 15.185 114.785 ;
        RECT 15.355 114.415 15.875 114.955 ;
        RECT 16.045 114.955 17.255 116.045 ;
        RECT 17.425 114.955 20.935 116.045 ;
        RECT 21.195 115.115 21.365 115.875 ;
        RECT 21.545 115.285 21.875 116.045 ;
        RECT 16.045 114.415 16.565 114.955 ;
        RECT 16.735 114.245 17.255 114.785 ;
        RECT 17.425 114.435 19.115 114.955 ;
        RECT 21.195 114.945 21.860 115.115 ;
        RECT 22.045 114.970 22.315 115.875 ;
        RECT 21.690 114.800 21.860 114.945 ;
        RECT 19.285 114.265 20.935 114.785 ;
        RECT 21.125 114.395 21.455 114.765 ;
        RECT 21.690 114.470 21.975 114.800 ;
        RECT 14.665 113.495 15.875 114.245 ;
        RECT 16.045 113.495 17.255 114.245 ;
        RECT 17.425 113.495 20.935 114.265 ;
        RECT 21.690 114.215 21.860 114.470 ;
        RECT 21.195 114.045 21.860 114.215 ;
        RECT 22.145 114.170 22.315 114.970 ;
        RECT 22.545 114.905 22.755 116.045 ;
        RECT 22.925 114.895 23.255 115.875 ;
        RECT 23.425 114.905 23.655 116.045 ;
        RECT 21.195 113.665 21.365 114.045 ;
        RECT 21.545 113.495 21.875 113.875 ;
        RECT 22.055 113.665 22.315 114.170 ;
        RECT 22.545 113.495 22.755 114.315 ;
        RECT 22.925 114.295 23.175 114.895 ;
        RECT 24.325 114.880 24.615 116.045 ;
        RECT 24.875 115.375 25.045 115.875 ;
        RECT 25.215 115.545 25.545 116.045 ;
        RECT 24.875 115.205 25.540 115.375 ;
        RECT 23.345 114.485 23.675 114.735 ;
        RECT 24.790 114.385 25.140 115.035 ;
        RECT 22.925 113.665 23.255 114.295 ;
        RECT 23.425 113.495 23.655 114.315 ;
        RECT 24.325 113.495 24.615 114.220 ;
        RECT 25.310 114.215 25.540 115.205 ;
        RECT 24.875 114.045 25.540 114.215 ;
        RECT 24.875 113.755 25.045 114.045 ;
        RECT 25.215 113.495 25.545 113.875 ;
        RECT 25.715 113.755 25.940 115.875 ;
        RECT 26.155 115.545 26.485 116.045 ;
        RECT 26.655 115.375 26.825 115.875 ;
        RECT 27.060 115.660 27.890 115.830 ;
        RECT 28.130 115.665 28.510 116.045 ;
        RECT 26.130 115.205 26.825 115.375 ;
        RECT 26.130 114.235 26.300 115.205 ;
        RECT 26.470 114.415 26.880 115.035 ;
        RECT 27.050 114.985 27.550 115.365 ;
        RECT 26.130 114.045 26.825 114.235 ;
        RECT 27.050 114.115 27.270 114.985 ;
        RECT 27.720 114.815 27.890 115.660 ;
        RECT 28.690 115.495 28.860 115.785 ;
        RECT 29.030 115.665 29.360 116.045 ;
        RECT 29.830 115.575 30.460 115.825 ;
        RECT 30.640 115.665 31.060 116.045 ;
        RECT 30.290 115.495 30.460 115.575 ;
        RECT 31.260 115.495 31.500 115.785 ;
        RECT 28.060 115.245 29.430 115.495 ;
        RECT 28.060 114.985 28.310 115.245 ;
        RECT 28.820 114.815 29.070 114.975 ;
        RECT 27.720 114.645 29.070 114.815 ;
        RECT 27.720 114.605 28.140 114.645 ;
        RECT 27.450 114.055 27.800 114.425 ;
        RECT 26.155 113.495 26.485 113.875 ;
        RECT 26.655 113.715 26.825 114.045 ;
        RECT 27.970 113.875 28.140 114.605 ;
        RECT 29.240 114.475 29.430 115.245 ;
        RECT 28.310 114.145 28.720 114.475 ;
        RECT 29.010 114.135 29.430 114.475 ;
        RECT 29.600 115.065 30.120 115.375 ;
        RECT 30.290 115.325 31.500 115.495 ;
        RECT 31.730 115.355 32.060 116.045 ;
        RECT 29.600 114.305 29.770 115.065 ;
        RECT 29.940 114.475 30.120 114.885 ;
        RECT 30.290 114.815 30.460 115.325 ;
        RECT 32.230 115.175 32.400 115.785 ;
        RECT 32.670 115.325 33.000 115.835 ;
        RECT 32.230 115.155 32.550 115.175 ;
        RECT 30.630 114.985 32.550 115.155 ;
        RECT 30.290 114.645 32.190 114.815 ;
        RECT 30.520 114.305 30.850 114.425 ;
        RECT 29.600 114.135 30.850 114.305 ;
        RECT 27.125 113.675 28.140 113.875 ;
        RECT 28.310 113.495 28.720 113.935 ;
        RECT 29.010 113.705 29.260 114.135 ;
        RECT 29.460 113.495 29.780 113.955 ;
        RECT 31.020 113.885 31.190 114.645 ;
        RECT 31.860 114.585 32.190 114.645 ;
        RECT 31.380 114.415 31.710 114.475 ;
        RECT 31.380 114.145 32.040 114.415 ;
        RECT 32.360 114.090 32.550 114.985 ;
        RECT 30.340 113.715 31.190 113.885 ;
        RECT 31.390 113.495 32.050 113.975 ;
        RECT 32.230 113.760 32.550 114.090 ;
        RECT 32.750 114.735 33.000 115.325 ;
        RECT 33.180 115.245 33.465 116.045 ;
        RECT 33.645 115.705 33.900 115.735 ;
        RECT 33.645 115.535 33.985 115.705 ;
        RECT 33.645 115.065 33.900 115.535 ;
        RECT 32.750 114.405 33.550 114.735 ;
        RECT 32.750 113.755 33.000 114.405 ;
        RECT 33.720 114.205 33.900 115.065 ;
        RECT 34.965 114.905 35.175 116.045 ;
        RECT 35.345 114.895 35.675 115.875 ;
        RECT 35.845 114.905 36.075 116.045 ;
        RECT 36.835 115.115 37.005 115.875 ;
        RECT 37.185 115.285 37.515 116.045 ;
        RECT 36.835 114.945 37.500 115.115 ;
        RECT 37.685 114.970 37.955 115.875 ;
        RECT 33.180 113.495 33.465 113.955 ;
        RECT 33.645 113.675 33.900 114.205 ;
        RECT 34.965 113.495 35.175 114.315 ;
        RECT 35.345 114.295 35.595 114.895 ;
        RECT 37.330 114.800 37.500 114.945 ;
        RECT 35.765 114.485 36.095 114.735 ;
        RECT 36.765 114.395 37.095 114.765 ;
        RECT 37.330 114.470 37.615 114.800 ;
        RECT 35.345 113.665 35.675 114.295 ;
        RECT 35.845 113.495 36.075 114.315 ;
        RECT 37.330 114.215 37.500 114.470 ;
        RECT 36.835 114.045 37.500 114.215 ;
        RECT 37.785 114.170 37.955 114.970 ;
        RECT 36.835 113.665 37.005 114.045 ;
        RECT 37.185 113.495 37.515 113.875 ;
        RECT 37.695 113.665 37.955 114.170 ;
        RECT 39.045 114.970 39.315 115.875 ;
        RECT 39.485 115.285 39.815 116.045 ;
        RECT 39.995 115.115 40.165 115.875 ;
        RECT 39.045 114.170 39.215 114.970 ;
        RECT 39.500 114.945 40.165 115.115 ;
        RECT 40.425 114.955 43.935 116.045 ;
        RECT 39.500 114.800 39.670 114.945 ;
        RECT 39.385 114.470 39.670 114.800 ;
        RECT 39.500 114.215 39.670 114.470 ;
        RECT 39.905 114.395 40.235 114.765 ;
        RECT 40.425 114.435 42.115 114.955 ;
        RECT 44.165 114.905 44.375 116.045 ;
        RECT 44.545 114.895 44.875 115.875 ;
        RECT 45.045 114.905 45.275 116.045 ;
        RECT 45.490 114.905 45.825 115.875 ;
        RECT 45.995 114.905 46.165 116.045 ;
        RECT 46.335 115.705 48.365 115.875 ;
        RECT 42.285 114.265 43.935 114.785 ;
        RECT 39.045 113.665 39.305 114.170 ;
        RECT 39.500 114.045 40.165 114.215 ;
        RECT 39.485 113.495 39.815 113.875 ;
        RECT 39.995 113.665 40.165 114.045 ;
        RECT 40.425 113.495 43.935 114.265 ;
        RECT 44.165 113.495 44.375 114.315 ;
        RECT 44.545 114.295 44.795 114.895 ;
        RECT 44.965 114.485 45.295 114.735 ;
        RECT 44.545 113.665 44.875 114.295 ;
        RECT 45.045 113.495 45.275 114.315 ;
        RECT 45.490 114.235 45.660 114.905 ;
        RECT 46.335 114.735 46.505 115.705 ;
        RECT 45.830 114.405 46.085 114.735 ;
        RECT 46.310 114.405 46.505 114.735 ;
        RECT 46.675 115.365 47.800 115.535 ;
        RECT 45.915 114.235 46.085 114.405 ;
        RECT 46.675 114.235 46.845 115.365 ;
        RECT 45.490 113.665 45.745 114.235 ;
        RECT 45.915 114.065 46.845 114.235 ;
        RECT 47.015 115.025 48.025 115.195 ;
        RECT 47.015 114.225 47.185 115.025 ;
        RECT 47.390 114.345 47.665 114.825 ;
        RECT 47.385 114.175 47.665 114.345 ;
        RECT 46.670 114.030 46.845 114.065 ;
        RECT 45.915 113.495 46.245 113.895 ;
        RECT 46.670 113.665 47.200 114.030 ;
        RECT 47.390 113.665 47.665 114.175 ;
        RECT 47.835 113.665 48.025 115.025 ;
        RECT 48.195 115.040 48.365 115.705 ;
        RECT 48.535 115.285 48.705 116.045 ;
        RECT 48.940 115.285 49.455 115.695 ;
        RECT 48.195 114.850 48.945 115.040 ;
        RECT 49.115 114.475 49.455 115.285 ;
        RECT 50.085 114.880 50.375 116.045 ;
        RECT 50.545 114.955 52.215 116.045 ;
        RECT 52.475 115.115 52.645 115.875 ;
        RECT 52.825 115.285 53.155 116.045 ;
        RECT 48.225 114.305 49.455 114.475 ;
        RECT 50.545 114.435 51.295 114.955 ;
        RECT 52.475 114.945 53.140 115.115 ;
        RECT 53.325 114.970 53.595 115.875 ;
        RECT 52.970 114.800 53.140 114.945 ;
        RECT 48.205 113.495 48.715 114.030 ;
        RECT 48.935 113.700 49.180 114.305 ;
        RECT 51.465 114.265 52.215 114.785 ;
        RECT 52.405 114.395 52.735 114.765 ;
        RECT 52.970 114.470 53.255 114.800 ;
        RECT 50.085 113.495 50.375 114.220 ;
        RECT 50.545 113.495 52.215 114.265 ;
        RECT 52.970 114.215 53.140 114.470 ;
        RECT 52.475 114.045 53.140 114.215 ;
        RECT 53.425 114.170 53.595 114.970 ;
        RECT 53.765 114.955 54.975 116.045 ;
        RECT 55.150 115.610 60.495 116.045 ;
        RECT 60.670 115.610 66.015 116.045 ;
        RECT 53.765 114.415 54.285 114.955 ;
        RECT 54.455 114.245 54.975 114.785 ;
        RECT 56.740 114.360 57.090 115.610 ;
        RECT 52.475 113.665 52.645 114.045 ;
        RECT 52.825 113.495 53.155 113.875 ;
        RECT 53.335 113.665 53.595 114.170 ;
        RECT 53.765 113.495 54.975 114.245 ;
        RECT 58.570 114.040 58.910 114.870 ;
        RECT 62.260 114.360 62.610 115.610 ;
        RECT 66.225 114.905 66.455 116.045 ;
        RECT 66.625 114.895 66.955 115.875 ;
        RECT 67.125 114.905 67.335 116.045 ;
        RECT 68.115 115.115 68.285 115.875 ;
        RECT 68.465 115.285 68.795 116.045 ;
        RECT 68.115 114.945 68.780 115.115 ;
        RECT 68.965 114.970 69.235 115.875 ;
        RECT 70.330 115.610 75.675 116.045 ;
        RECT 64.090 114.040 64.430 114.870 ;
        RECT 66.205 114.485 66.535 114.735 ;
        RECT 55.150 113.495 60.495 114.040 ;
        RECT 60.670 113.495 66.015 114.040 ;
        RECT 66.225 113.495 66.455 114.315 ;
        RECT 66.705 114.295 66.955 114.895 ;
        RECT 68.610 114.800 68.780 114.945 ;
        RECT 68.045 114.395 68.375 114.765 ;
        RECT 68.610 114.470 68.895 114.800 ;
        RECT 66.625 113.665 66.955 114.295 ;
        RECT 67.125 113.495 67.335 114.315 ;
        RECT 68.610 114.215 68.780 114.470 ;
        RECT 68.115 114.045 68.780 114.215 ;
        RECT 69.065 114.170 69.235 114.970 ;
        RECT 71.920 114.360 72.270 115.610 ;
        RECT 75.845 114.880 76.135 116.045 ;
        RECT 77.600 115.705 77.855 115.735 ;
        RECT 77.515 115.535 77.855 115.705 ;
        RECT 77.600 115.065 77.855 115.535 ;
        RECT 78.035 115.245 78.320 116.045 ;
        RECT 78.500 115.325 78.830 115.835 ;
        RECT 68.115 113.665 68.285 114.045 ;
        RECT 68.465 113.495 68.795 113.875 ;
        RECT 68.975 113.665 69.235 114.170 ;
        RECT 73.750 114.040 74.090 114.870 ;
        RECT 70.330 113.495 75.675 114.040 ;
        RECT 75.845 113.495 76.135 114.220 ;
        RECT 77.600 114.205 77.780 115.065 ;
        RECT 78.500 114.735 78.750 115.325 ;
        RECT 79.100 115.175 79.270 115.785 ;
        RECT 79.440 115.355 79.770 116.045 ;
        RECT 80.000 115.495 80.240 115.785 ;
        RECT 80.440 115.665 80.860 116.045 ;
        RECT 81.040 115.575 81.670 115.825 ;
        RECT 82.140 115.665 82.470 116.045 ;
        RECT 81.040 115.495 81.210 115.575 ;
        RECT 82.640 115.495 82.810 115.785 ;
        RECT 82.990 115.665 83.370 116.045 ;
        RECT 83.610 115.660 84.440 115.830 ;
        RECT 80.000 115.325 81.210 115.495 ;
        RECT 77.950 114.405 78.750 114.735 ;
        RECT 77.600 113.675 77.855 114.205 ;
        RECT 78.035 113.495 78.320 113.955 ;
        RECT 78.500 113.755 78.750 114.405 ;
        RECT 78.950 115.155 79.270 115.175 ;
        RECT 78.950 114.985 80.870 115.155 ;
        RECT 78.950 114.090 79.140 114.985 ;
        RECT 81.040 114.815 81.210 115.325 ;
        RECT 81.380 115.065 81.900 115.375 ;
        RECT 79.310 114.645 81.210 114.815 ;
        RECT 79.310 114.585 79.640 114.645 ;
        RECT 79.790 114.415 80.120 114.475 ;
        RECT 79.460 114.145 80.120 114.415 ;
        RECT 78.950 113.760 79.270 114.090 ;
        RECT 79.450 113.495 80.110 113.975 ;
        RECT 80.310 113.885 80.480 114.645 ;
        RECT 81.380 114.475 81.560 114.885 ;
        RECT 80.650 114.305 80.980 114.425 ;
        RECT 81.730 114.305 81.900 115.065 ;
        RECT 80.650 114.135 81.900 114.305 ;
        RECT 82.070 115.245 83.440 115.495 ;
        RECT 82.070 114.475 82.260 115.245 ;
        RECT 83.190 114.985 83.440 115.245 ;
        RECT 82.430 114.815 82.680 114.975 ;
        RECT 83.610 114.815 83.780 115.660 ;
        RECT 84.675 115.375 84.845 115.875 ;
        RECT 85.015 115.545 85.345 116.045 ;
        RECT 83.950 114.985 84.450 115.365 ;
        RECT 84.675 115.205 85.370 115.375 ;
        RECT 82.430 114.645 83.780 114.815 ;
        RECT 83.360 114.605 83.780 114.645 ;
        RECT 82.070 114.135 82.490 114.475 ;
        RECT 82.780 114.145 83.190 114.475 ;
        RECT 80.310 113.715 81.160 113.885 ;
        RECT 81.720 113.495 82.040 113.955 ;
        RECT 82.240 113.705 82.490 114.135 ;
        RECT 82.780 113.495 83.190 113.935 ;
        RECT 83.360 113.875 83.530 114.605 ;
        RECT 83.700 114.055 84.050 114.425 ;
        RECT 84.230 114.115 84.450 114.985 ;
        RECT 84.620 114.415 85.030 115.035 ;
        RECT 85.200 114.235 85.370 115.205 ;
        RECT 84.675 114.045 85.370 114.235 ;
        RECT 83.360 113.675 84.375 113.875 ;
        RECT 84.675 113.715 84.845 114.045 ;
        RECT 85.015 113.495 85.345 113.875 ;
        RECT 85.560 113.755 85.785 115.875 ;
        RECT 85.955 115.545 86.285 116.045 ;
        RECT 86.455 115.375 86.625 115.875 ;
        RECT 85.960 115.205 86.625 115.375 ;
        RECT 87.435 115.375 87.605 115.875 ;
        RECT 87.775 115.545 88.105 116.045 ;
        RECT 87.435 115.205 88.100 115.375 ;
        RECT 85.960 114.215 86.190 115.205 ;
        RECT 86.360 114.385 86.710 115.035 ;
        RECT 87.350 114.385 87.700 115.035 ;
        RECT 87.870 114.215 88.100 115.205 ;
        RECT 85.960 114.045 86.625 114.215 ;
        RECT 85.955 113.495 86.285 113.875 ;
        RECT 86.455 113.755 86.625 114.045 ;
        RECT 87.435 114.045 88.100 114.215 ;
        RECT 87.435 113.755 87.605 114.045 ;
        RECT 87.775 113.495 88.105 113.875 ;
        RECT 88.275 113.755 88.500 115.875 ;
        RECT 88.715 115.545 89.045 116.045 ;
        RECT 89.215 115.375 89.385 115.875 ;
        RECT 89.620 115.660 90.450 115.830 ;
        RECT 90.690 115.665 91.070 116.045 ;
        RECT 88.690 115.205 89.385 115.375 ;
        RECT 88.690 114.235 88.860 115.205 ;
        RECT 89.030 114.415 89.440 115.035 ;
        RECT 89.610 114.985 90.110 115.365 ;
        RECT 88.690 114.045 89.385 114.235 ;
        RECT 89.610 114.115 89.830 114.985 ;
        RECT 90.280 114.815 90.450 115.660 ;
        RECT 91.250 115.495 91.420 115.785 ;
        RECT 91.590 115.665 91.920 116.045 ;
        RECT 92.390 115.575 93.020 115.825 ;
        RECT 93.200 115.665 93.620 116.045 ;
        RECT 92.850 115.495 93.020 115.575 ;
        RECT 93.820 115.495 94.060 115.785 ;
        RECT 90.620 115.245 91.990 115.495 ;
        RECT 90.620 114.985 90.870 115.245 ;
        RECT 91.380 114.815 91.630 114.975 ;
        RECT 90.280 114.645 91.630 114.815 ;
        RECT 90.280 114.605 90.700 114.645 ;
        RECT 90.010 114.055 90.360 114.425 ;
        RECT 88.715 113.495 89.045 113.875 ;
        RECT 89.215 113.715 89.385 114.045 ;
        RECT 90.530 113.875 90.700 114.605 ;
        RECT 91.800 114.475 91.990 115.245 ;
        RECT 90.870 114.145 91.280 114.475 ;
        RECT 91.570 114.135 91.990 114.475 ;
        RECT 92.160 115.065 92.680 115.375 ;
        RECT 92.850 115.325 94.060 115.495 ;
        RECT 94.290 115.355 94.620 116.045 ;
        RECT 92.160 114.305 92.330 115.065 ;
        RECT 92.500 114.475 92.680 114.885 ;
        RECT 92.850 114.815 93.020 115.325 ;
        RECT 94.790 115.175 94.960 115.785 ;
        RECT 95.230 115.325 95.560 115.835 ;
        RECT 94.790 115.155 95.110 115.175 ;
        RECT 93.190 114.985 95.110 115.155 ;
        RECT 92.850 114.645 94.750 114.815 ;
        RECT 93.080 114.305 93.410 114.425 ;
        RECT 92.160 114.135 93.410 114.305 ;
        RECT 89.685 113.675 90.700 113.875 ;
        RECT 90.870 113.495 91.280 113.935 ;
        RECT 91.570 113.705 91.820 114.135 ;
        RECT 92.020 113.495 92.340 113.955 ;
        RECT 93.580 113.885 93.750 114.645 ;
        RECT 94.420 114.585 94.750 114.645 ;
        RECT 93.940 114.415 94.270 114.475 ;
        RECT 93.940 114.145 94.600 114.415 ;
        RECT 94.920 114.090 95.110 114.985 ;
        RECT 92.900 113.715 93.750 113.885 ;
        RECT 93.950 113.495 94.610 113.975 ;
        RECT 94.790 113.760 95.110 114.090 ;
        RECT 95.310 114.735 95.560 115.325 ;
        RECT 95.740 115.245 96.025 116.045 ;
        RECT 96.205 115.705 96.460 115.735 ;
        RECT 96.205 115.535 96.545 115.705 ;
        RECT 96.205 115.065 96.460 115.535 ;
        RECT 95.310 114.405 96.110 114.735 ;
        RECT 95.310 113.755 95.560 114.405 ;
        RECT 96.280 114.205 96.460 115.065 ;
        RECT 97.465 114.955 100.055 116.045 ;
        RECT 100.225 114.970 100.495 115.875 ;
        RECT 100.665 115.285 100.995 116.045 ;
        RECT 101.175 115.115 101.345 115.875 ;
        RECT 97.465 114.435 98.675 114.955 ;
        RECT 98.845 114.265 100.055 114.785 ;
        RECT 95.740 113.495 96.025 113.955 ;
        RECT 96.205 113.675 96.460 114.205 ;
        RECT 97.465 113.495 100.055 114.265 ;
        RECT 100.225 114.170 100.395 114.970 ;
        RECT 100.680 114.945 101.345 115.115 ;
        RECT 100.680 114.800 100.850 114.945 ;
        RECT 101.605 114.880 101.895 116.045 ;
        RECT 102.530 115.610 107.875 116.045 ;
        RECT 100.565 114.470 100.850 114.800 ;
        RECT 100.680 114.215 100.850 114.470 ;
        RECT 101.085 114.395 101.415 114.765 ;
        RECT 104.120 114.360 104.470 115.610 ;
        RECT 108.135 115.115 108.305 115.875 ;
        RECT 108.485 115.285 108.815 116.045 ;
        RECT 108.135 114.945 108.800 115.115 ;
        RECT 108.985 114.970 109.255 115.875 ;
        RECT 100.225 113.665 100.485 114.170 ;
        RECT 100.680 114.045 101.345 114.215 ;
        RECT 100.665 113.495 100.995 113.875 ;
        RECT 101.175 113.665 101.345 114.045 ;
        RECT 101.605 113.495 101.895 114.220 ;
        RECT 105.950 114.040 106.290 114.870 ;
        RECT 108.630 114.800 108.800 114.945 ;
        RECT 108.065 114.395 108.395 114.765 ;
        RECT 108.630 114.470 108.915 114.800 ;
        RECT 108.630 114.215 108.800 114.470 ;
        RECT 108.135 114.045 108.800 114.215 ;
        RECT 109.085 114.170 109.255 114.970 ;
        RECT 109.425 114.955 111.095 116.045 ;
        RECT 111.265 115.285 111.780 115.695 ;
        RECT 112.015 115.285 112.185 116.045 ;
        RECT 112.355 115.705 114.385 115.875 ;
        RECT 109.425 114.435 110.175 114.955 ;
        RECT 110.345 114.265 111.095 114.785 ;
        RECT 111.265 114.475 111.605 115.285 ;
        RECT 112.355 115.040 112.525 115.705 ;
        RECT 112.920 115.365 114.045 115.535 ;
        RECT 111.775 114.850 112.525 115.040 ;
        RECT 112.695 115.025 113.705 115.195 ;
        RECT 111.265 114.305 112.495 114.475 ;
        RECT 102.530 113.495 107.875 114.040 ;
        RECT 108.135 113.665 108.305 114.045 ;
        RECT 108.485 113.495 108.815 113.875 ;
        RECT 108.995 113.665 109.255 114.170 ;
        RECT 109.425 113.495 111.095 114.265 ;
        RECT 111.540 113.700 111.785 114.305 ;
        RECT 112.005 113.495 112.515 114.030 ;
        RECT 112.695 113.665 112.885 115.025 ;
        RECT 113.055 114.685 113.330 114.825 ;
        RECT 113.055 114.515 113.335 114.685 ;
        RECT 113.055 113.665 113.330 114.515 ;
        RECT 113.535 114.225 113.705 115.025 ;
        RECT 113.875 114.235 114.045 115.365 ;
        RECT 114.215 114.735 114.385 115.705 ;
        RECT 114.555 114.905 114.725 116.045 ;
        RECT 114.895 114.905 115.230 115.875 ;
        RECT 115.410 115.610 120.755 116.045 ;
        RECT 120.930 115.610 126.275 116.045 ;
        RECT 114.215 114.405 114.410 114.735 ;
        RECT 114.635 114.405 114.890 114.735 ;
        RECT 114.635 114.235 114.805 114.405 ;
        RECT 115.060 114.235 115.230 114.905 ;
        RECT 117.000 114.360 117.350 115.610 ;
        RECT 113.875 114.065 114.805 114.235 ;
        RECT 113.875 114.030 114.050 114.065 ;
        RECT 113.520 113.665 114.050 114.030 ;
        RECT 114.475 113.495 114.805 113.895 ;
        RECT 114.975 113.665 115.230 114.235 ;
        RECT 118.830 114.040 119.170 114.870 ;
        RECT 122.520 114.360 122.870 115.610 ;
        RECT 126.445 114.955 127.655 116.045 ;
        RECT 124.350 114.040 124.690 114.870 ;
        RECT 126.445 114.415 126.965 114.955 ;
        RECT 127.135 114.245 127.655 114.785 ;
        RECT 115.410 113.495 120.755 114.040 ;
        RECT 120.930 113.495 126.275 114.040 ;
        RECT 126.445 113.495 127.655 114.245 ;
        RECT 14.580 113.325 127.740 113.495 ;
        RECT 14.665 112.575 15.875 113.325 ;
        RECT 16.355 112.855 16.525 113.325 ;
        RECT 16.695 112.675 17.025 113.155 ;
        RECT 17.195 112.855 17.365 113.325 ;
        RECT 17.535 112.675 17.865 113.155 ;
        RECT 14.665 112.035 15.185 112.575 ;
        RECT 16.100 112.505 17.865 112.675 ;
        RECT 18.035 112.515 18.205 113.325 ;
        RECT 18.405 112.945 19.475 113.115 ;
        RECT 18.405 112.590 18.725 112.945 ;
        RECT 15.355 111.865 15.875 112.405 ;
        RECT 14.665 110.775 15.875 111.865 ;
        RECT 16.100 111.955 16.510 112.505 ;
        RECT 18.400 112.335 18.725 112.590 ;
        RECT 16.695 112.125 18.725 112.335 ;
        RECT 18.380 112.115 18.725 112.125 ;
        RECT 18.895 112.375 19.135 112.775 ;
        RECT 19.305 112.715 19.475 112.945 ;
        RECT 19.645 112.885 19.835 113.325 ;
        RECT 20.005 112.875 20.955 113.155 ;
        RECT 21.175 112.965 21.525 113.135 ;
        RECT 19.305 112.545 19.835 112.715 ;
        RECT 16.100 111.785 17.825 111.955 ;
        RECT 16.355 110.775 16.525 111.615 ;
        RECT 16.735 110.945 16.985 111.785 ;
        RECT 17.195 110.775 17.365 111.615 ;
        RECT 17.535 110.945 17.825 111.785 ;
        RECT 18.035 110.775 18.205 111.835 ;
        RECT 18.380 111.495 18.550 112.115 ;
        RECT 18.895 112.005 19.435 112.375 ;
        RECT 19.615 112.265 19.835 112.545 ;
        RECT 20.005 112.095 20.175 112.875 ;
        RECT 19.770 111.925 20.175 112.095 ;
        RECT 20.345 112.085 20.695 112.705 ;
        RECT 19.770 111.835 19.940 111.925 ;
        RECT 20.865 111.915 21.075 112.705 ;
        RECT 18.720 111.665 19.940 111.835 ;
        RECT 20.400 111.755 21.075 111.915 ;
        RECT 18.380 111.325 19.180 111.495 ;
        RECT 18.500 110.775 18.830 111.155 ;
        RECT 19.010 111.035 19.180 111.325 ;
        RECT 19.770 111.285 19.940 111.665 ;
        RECT 20.110 111.745 21.075 111.755 ;
        RECT 21.265 112.575 21.525 112.965 ;
        RECT 21.735 112.865 22.065 113.325 ;
        RECT 22.940 112.935 23.795 113.105 ;
        RECT 24.000 112.935 24.495 113.105 ;
        RECT 24.665 112.965 24.995 113.325 ;
        RECT 21.265 111.885 21.435 112.575 ;
        RECT 21.605 112.225 21.775 112.405 ;
        RECT 21.945 112.395 22.735 112.645 ;
        RECT 22.940 112.225 23.110 112.935 ;
        RECT 23.280 112.425 23.635 112.645 ;
        RECT 21.605 112.055 23.295 112.225 ;
        RECT 20.110 111.455 20.570 111.745 ;
        RECT 21.265 111.715 22.765 111.885 ;
        RECT 21.265 111.575 21.435 111.715 ;
        RECT 20.875 111.405 21.435 111.575 ;
        RECT 19.350 110.775 19.600 111.235 ;
        RECT 19.770 110.945 20.640 111.285 ;
        RECT 20.875 110.945 21.045 111.405 ;
        RECT 21.880 111.375 22.955 111.545 ;
        RECT 21.215 110.775 21.585 111.235 ;
        RECT 21.880 111.035 22.050 111.375 ;
        RECT 22.220 110.775 22.550 111.205 ;
        RECT 22.785 111.035 22.955 111.375 ;
        RECT 23.125 111.275 23.295 112.055 ;
        RECT 23.465 111.835 23.635 112.425 ;
        RECT 23.805 112.025 24.155 112.645 ;
        RECT 23.465 111.445 23.930 111.835 ;
        RECT 24.325 111.575 24.495 112.935 ;
        RECT 24.665 111.745 25.125 112.795 ;
        RECT 24.100 111.405 24.495 111.575 ;
        RECT 24.100 111.275 24.270 111.405 ;
        RECT 23.125 110.945 23.805 111.275 ;
        RECT 24.020 110.945 24.270 111.275 ;
        RECT 24.440 110.775 24.690 111.235 ;
        RECT 24.860 110.960 25.185 111.745 ;
        RECT 25.355 110.945 25.525 113.065 ;
        RECT 25.695 112.945 26.025 113.325 ;
        RECT 26.195 112.775 26.450 113.065 ;
        RECT 25.700 112.605 26.450 112.775 ;
        RECT 25.700 111.615 25.930 112.605 ;
        RECT 26.625 112.555 28.295 113.325 ;
        RECT 28.470 112.780 33.815 113.325 ;
        RECT 26.100 111.785 26.450 112.435 ;
        RECT 26.625 111.865 27.375 112.385 ;
        RECT 27.545 112.035 28.295 112.555 ;
        RECT 25.700 111.445 26.450 111.615 ;
        RECT 25.695 110.775 26.025 111.275 ;
        RECT 26.195 110.945 26.450 111.445 ;
        RECT 26.625 110.775 28.295 111.865 ;
        RECT 30.060 111.210 30.410 112.460 ;
        RECT 31.890 111.950 32.230 112.780 ;
        RECT 34.045 112.505 34.255 113.325 ;
        RECT 34.425 112.525 34.755 113.155 ;
        RECT 34.425 111.925 34.675 112.525 ;
        RECT 34.925 112.505 35.155 113.325 ;
        RECT 35.365 112.555 37.035 113.325 ;
        RECT 37.205 112.600 37.495 113.325 ;
        RECT 38.215 112.845 38.515 113.325 ;
        RECT 38.685 112.675 38.945 113.130 ;
        RECT 39.115 112.845 39.375 113.325 ;
        RECT 39.555 112.675 39.815 113.130 ;
        RECT 39.985 112.845 40.235 113.325 ;
        RECT 40.415 112.675 40.675 113.130 ;
        RECT 40.845 112.845 41.095 113.325 ;
        RECT 41.275 112.675 41.535 113.130 ;
        RECT 41.705 112.845 41.950 113.325 ;
        RECT 42.120 112.675 42.395 113.130 ;
        RECT 42.565 112.845 42.810 113.325 ;
        RECT 42.980 112.675 43.240 113.130 ;
        RECT 43.410 112.845 43.670 113.325 ;
        RECT 43.840 112.675 44.100 113.130 ;
        RECT 44.270 112.845 44.530 113.325 ;
        RECT 44.700 112.675 44.960 113.130 ;
        RECT 45.130 112.765 45.390 113.325 ;
        RECT 34.845 112.085 35.175 112.335 ;
        RECT 28.470 110.775 33.815 111.210 ;
        RECT 34.045 110.775 34.255 111.915 ;
        RECT 34.425 110.945 34.755 111.925 ;
        RECT 34.925 110.775 35.155 111.915 ;
        RECT 35.365 111.865 36.115 112.385 ;
        RECT 36.285 112.035 37.035 112.555 ;
        RECT 38.215 112.505 44.960 112.675 ;
        RECT 35.365 110.775 37.035 111.865 ;
        RECT 37.205 110.775 37.495 111.940 ;
        RECT 38.215 111.915 39.380 112.505 ;
        RECT 45.560 112.335 45.810 113.145 ;
        RECT 45.990 112.800 46.250 113.325 ;
        RECT 46.420 112.335 46.670 113.145 ;
        RECT 46.850 112.815 47.155 113.325 ;
        RECT 39.550 112.085 46.670 112.335 ;
        RECT 46.840 112.085 47.155 112.645 ;
        RECT 48.245 112.555 51.755 113.325 ;
        RECT 51.930 112.780 57.275 113.325 ;
        RECT 57.450 112.780 62.795 113.325 ;
        RECT 38.215 111.690 44.960 111.915 ;
        RECT 38.215 110.775 38.485 111.520 ;
        RECT 38.655 110.950 38.945 111.690 ;
        RECT 39.555 111.675 44.960 111.690 ;
        RECT 39.115 110.780 39.370 111.505 ;
        RECT 39.555 110.950 39.815 111.675 ;
        RECT 39.985 110.780 40.230 111.505 ;
        RECT 40.415 110.950 40.675 111.675 ;
        RECT 40.845 110.780 41.090 111.505 ;
        RECT 41.275 110.950 41.535 111.675 ;
        RECT 41.705 110.780 41.950 111.505 ;
        RECT 42.120 110.950 42.380 111.675 ;
        RECT 42.550 110.780 42.810 111.505 ;
        RECT 42.980 110.950 43.240 111.675 ;
        RECT 43.410 110.780 43.670 111.505 ;
        RECT 43.840 110.950 44.100 111.675 ;
        RECT 44.270 110.780 44.530 111.505 ;
        RECT 44.700 110.950 44.960 111.675 ;
        RECT 45.130 110.780 45.390 111.575 ;
        RECT 45.560 110.950 45.810 112.085 ;
        RECT 39.115 110.775 45.390 110.780 ;
        RECT 45.990 110.775 46.250 111.585 ;
        RECT 46.425 110.945 46.670 112.085 ;
        RECT 48.245 111.865 49.935 112.385 ;
        RECT 50.105 112.035 51.755 112.555 ;
        RECT 46.850 110.775 47.145 111.585 ;
        RECT 48.245 110.775 51.755 111.865 ;
        RECT 53.520 111.210 53.870 112.460 ;
        RECT 55.350 111.950 55.690 112.780 ;
        RECT 59.040 111.210 59.390 112.460 ;
        RECT 60.870 111.950 61.210 112.780 ;
        RECT 62.965 112.600 63.255 113.325 ;
        RECT 63.890 112.780 69.235 113.325 ;
        RECT 69.410 112.780 74.755 113.325 ;
        RECT 74.930 112.780 80.275 113.325 ;
        RECT 51.930 110.775 57.275 111.210 ;
        RECT 57.450 110.775 62.795 111.210 ;
        RECT 62.965 110.775 63.255 111.940 ;
        RECT 65.480 111.210 65.830 112.460 ;
        RECT 67.310 111.950 67.650 112.780 ;
        RECT 71.000 111.210 71.350 112.460 ;
        RECT 72.830 111.950 73.170 112.780 ;
        RECT 76.520 111.210 76.870 112.460 ;
        RECT 78.350 111.950 78.690 112.780 ;
        RECT 80.505 112.505 80.715 113.325 ;
        RECT 80.885 112.525 81.215 113.155 ;
        RECT 80.885 111.925 81.135 112.525 ;
        RECT 81.385 112.505 81.615 113.325 ;
        RECT 81.825 112.575 83.035 113.325 ;
        RECT 83.210 112.780 88.555 113.325 ;
        RECT 81.305 112.085 81.635 112.335 ;
        RECT 63.890 110.775 69.235 111.210 ;
        RECT 69.410 110.775 74.755 111.210 ;
        RECT 74.930 110.775 80.275 111.210 ;
        RECT 80.505 110.775 80.715 111.915 ;
        RECT 80.885 110.945 81.215 111.925 ;
        RECT 81.385 110.775 81.615 111.915 ;
        RECT 81.825 111.865 82.345 112.405 ;
        RECT 82.515 112.035 83.035 112.575 ;
        RECT 81.825 110.775 83.035 111.865 ;
        RECT 84.800 111.210 85.150 112.460 ;
        RECT 86.630 111.950 86.970 112.780 ;
        RECT 88.725 112.600 89.015 113.325 ;
        RECT 89.185 112.555 92.695 113.325 ;
        RECT 92.865 112.815 93.170 113.325 ;
        RECT 83.210 110.775 88.555 111.210 ;
        RECT 88.725 110.775 89.015 111.940 ;
        RECT 89.185 111.865 90.875 112.385 ;
        RECT 91.045 112.035 92.695 112.555 ;
        RECT 92.865 112.085 93.180 112.645 ;
        RECT 93.350 112.335 93.600 113.145 ;
        RECT 93.770 112.800 94.030 113.325 ;
        RECT 94.210 112.335 94.460 113.145 ;
        RECT 94.630 112.765 94.890 113.325 ;
        RECT 95.060 112.675 95.320 113.130 ;
        RECT 95.490 112.845 95.750 113.325 ;
        RECT 95.920 112.675 96.180 113.130 ;
        RECT 96.350 112.845 96.610 113.325 ;
        RECT 96.780 112.675 97.040 113.130 ;
        RECT 97.210 112.845 97.455 113.325 ;
        RECT 97.625 112.675 97.900 113.130 ;
        RECT 98.070 112.845 98.315 113.325 ;
        RECT 98.485 112.675 98.745 113.130 ;
        RECT 98.925 112.845 99.175 113.325 ;
        RECT 99.345 112.675 99.605 113.130 ;
        RECT 99.785 112.845 100.035 113.325 ;
        RECT 100.205 112.675 100.465 113.130 ;
        RECT 100.645 112.845 100.905 113.325 ;
        RECT 101.075 112.675 101.335 113.130 ;
        RECT 101.505 112.845 101.805 113.325 ;
        RECT 102.065 112.820 102.350 113.325 ;
        RECT 95.060 112.645 101.805 112.675 ;
        RECT 102.520 112.650 102.845 113.155 ;
        RECT 95.060 112.505 101.835 112.645 ;
        RECT 100.640 112.475 101.835 112.505 ;
        RECT 93.350 112.085 100.470 112.335 ;
        RECT 89.185 110.775 92.695 111.865 ;
        RECT 92.875 110.775 93.170 111.585 ;
        RECT 93.350 110.945 93.595 112.085 ;
        RECT 93.770 110.775 94.030 111.585 ;
        RECT 94.210 110.950 94.460 112.085 ;
        RECT 100.640 111.915 101.805 112.475 ;
        RECT 102.065 112.120 102.845 112.650 ;
        RECT 95.060 111.690 101.805 111.915 ;
        RECT 95.060 111.675 100.465 111.690 ;
        RECT 94.630 110.780 94.890 111.575 ;
        RECT 95.060 110.950 95.320 111.675 ;
        RECT 95.490 110.780 95.750 111.505 ;
        RECT 95.920 110.950 96.180 111.675 ;
        RECT 96.350 110.780 96.610 111.505 ;
        RECT 96.780 110.950 97.040 111.675 ;
        RECT 97.210 110.780 97.470 111.505 ;
        RECT 97.640 110.950 97.900 111.675 ;
        RECT 98.070 110.780 98.315 111.505 ;
        RECT 98.485 110.950 98.745 111.675 ;
        RECT 98.930 110.780 99.175 111.505 ;
        RECT 99.345 110.950 99.605 111.675 ;
        RECT 99.790 110.780 100.035 111.505 ;
        RECT 100.205 110.950 100.465 111.675 ;
        RECT 100.650 110.780 100.905 111.505 ;
        RECT 101.075 110.950 101.365 111.690 ;
        RECT 94.630 110.775 100.905 110.780 ;
        RECT 101.535 110.775 101.805 111.520 ;
        RECT 102.065 110.775 102.345 111.745 ;
        RECT 102.515 110.945 102.845 112.120 ;
        RECT 103.035 112.085 103.275 113.035 ;
        RECT 103.450 112.780 108.795 113.325 ;
        RECT 108.970 112.780 114.315 113.325 ;
        RECT 103.015 110.775 103.275 111.745 ;
        RECT 105.040 111.210 105.390 112.460 ;
        RECT 106.870 111.950 107.210 112.780 ;
        RECT 110.560 111.210 110.910 112.460 ;
        RECT 112.390 111.950 112.730 112.780 ;
        RECT 114.485 112.600 114.775 113.325 ;
        RECT 115.865 112.555 119.375 113.325 ;
        RECT 103.450 110.775 108.795 111.210 ;
        RECT 108.970 110.775 114.315 111.210 ;
        RECT 114.485 110.775 114.775 111.940 ;
        RECT 115.865 111.865 117.555 112.385 ;
        RECT 117.725 112.035 119.375 112.555 ;
        RECT 119.585 112.505 119.815 113.325 ;
        RECT 119.985 112.525 120.315 113.155 ;
        RECT 119.565 112.085 119.895 112.335 ;
        RECT 120.065 111.925 120.315 112.525 ;
        RECT 120.485 112.505 120.695 113.325 ;
        RECT 120.925 112.650 121.185 113.155 ;
        RECT 121.365 112.945 121.695 113.325 ;
        RECT 121.875 112.775 122.045 113.155 ;
        RECT 115.865 110.775 119.375 111.865 ;
        RECT 119.585 110.775 119.815 111.915 ;
        RECT 119.985 110.945 120.315 111.925 ;
        RECT 120.485 110.775 120.695 111.915 ;
        RECT 120.925 111.850 121.095 112.650 ;
        RECT 121.380 112.605 122.045 112.775 ;
        RECT 122.305 112.650 122.565 113.155 ;
        RECT 122.745 112.945 123.075 113.325 ;
        RECT 123.255 112.775 123.425 113.155 ;
        RECT 121.380 112.350 121.550 112.605 ;
        RECT 121.265 112.020 121.550 112.350 ;
        RECT 121.785 112.055 122.115 112.425 ;
        RECT 121.380 111.875 121.550 112.020 ;
        RECT 120.925 110.945 121.195 111.850 ;
        RECT 121.380 111.705 122.045 111.875 ;
        RECT 121.365 110.775 121.695 111.535 ;
        RECT 121.875 110.945 122.045 111.705 ;
        RECT 122.305 111.850 122.475 112.650 ;
        RECT 122.760 112.605 123.425 112.775 ;
        RECT 122.760 112.350 122.930 112.605 ;
        RECT 123.685 112.555 126.275 113.325 ;
        RECT 126.445 112.575 127.655 113.325 ;
        RECT 122.645 112.020 122.930 112.350 ;
        RECT 123.165 112.055 123.495 112.425 ;
        RECT 122.760 111.875 122.930 112.020 ;
        RECT 122.305 110.945 122.575 111.850 ;
        RECT 122.760 111.705 123.425 111.875 ;
        RECT 122.745 110.775 123.075 111.535 ;
        RECT 123.255 110.945 123.425 111.705 ;
        RECT 123.685 111.865 124.895 112.385 ;
        RECT 125.065 112.035 126.275 112.555 ;
        RECT 126.445 111.865 126.965 112.405 ;
        RECT 127.135 112.035 127.655 112.575 ;
        RECT 123.685 110.775 126.275 111.865 ;
        RECT 126.445 110.775 127.655 111.865 ;
        RECT 14.580 110.605 127.740 110.775 ;
        RECT 14.665 109.515 15.875 110.605 ;
        RECT 14.665 108.805 15.185 109.345 ;
        RECT 15.355 108.975 15.875 109.515 ;
        RECT 16.965 109.515 20.475 110.605 ;
        RECT 16.965 108.995 18.655 109.515 ;
        RECT 20.705 109.465 20.915 110.605 ;
        RECT 21.085 109.455 21.415 110.435 ;
        RECT 21.585 109.465 21.815 110.605 ;
        RECT 23.005 109.465 23.215 110.605 ;
        RECT 23.385 109.455 23.715 110.435 ;
        RECT 23.885 109.465 24.115 110.605 ;
        RECT 18.825 108.825 20.475 109.345 ;
        RECT 14.665 108.055 15.875 108.805 ;
        RECT 16.965 108.055 20.475 108.825 ;
        RECT 20.705 108.055 20.915 108.875 ;
        RECT 21.085 108.855 21.335 109.455 ;
        RECT 21.505 109.045 21.835 109.295 ;
        RECT 21.085 108.225 21.415 108.855 ;
        RECT 21.585 108.055 21.815 108.875 ;
        RECT 23.005 108.055 23.215 108.875 ;
        RECT 23.385 108.855 23.635 109.455 ;
        RECT 24.325 109.440 24.615 110.605 ;
        RECT 24.785 109.515 27.375 110.605 ;
        RECT 27.545 109.530 27.815 110.435 ;
        RECT 27.985 109.845 28.315 110.605 ;
        RECT 28.495 109.675 28.665 110.435 ;
        RECT 23.805 109.045 24.135 109.295 ;
        RECT 24.785 108.995 25.995 109.515 ;
        RECT 23.385 108.225 23.715 108.855 ;
        RECT 23.885 108.055 24.115 108.875 ;
        RECT 26.165 108.825 27.375 109.345 ;
        RECT 24.325 108.055 24.615 108.780 ;
        RECT 24.785 108.055 27.375 108.825 ;
        RECT 27.545 108.730 27.715 109.530 ;
        RECT 28.000 109.505 28.665 109.675 ;
        RECT 28.925 109.515 30.595 110.605 ;
        RECT 28.000 109.360 28.170 109.505 ;
        RECT 27.885 109.030 28.170 109.360 ;
        RECT 28.000 108.775 28.170 109.030 ;
        RECT 28.405 108.955 28.735 109.325 ;
        RECT 28.925 108.995 29.675 109.515 ;
        RECT 30.825 109.465 31.035 110.605 ;
        RECT 31.205 109.455 31.535 110.435 ;
        RECT 31.705 109.465 31.935 110.605 ;
        RECT 32.145 109.530 32.415 110.435 ;
        RECT 32.585 109.845 32.915 110.605 ;
        RECT 33.095 109.675 33.265 110.435 ;
        RECT 29.845 108.825 30.595 109.345 ;
        RECT 27.545 108.225 27.805 108.730 ;
        RECT 28.000 108.605 28.665 108.775 ;
        RECT 27.985 108.055 28.315 108.435 ;
        RECT 28.495 108.225 28.665 108.605 ;
        RECT 28.925 108.055 30.595 108.825 ;
        RECT 30.825 108.055 31.035 108.875 ;
        RECT 31.205 108.855 31.455 109.455 ;
        RECT 31.625 109.045 31.955 109.295 ;
        RECT 31.205 108.225 31.535 108.855 ;
        RECT 31.705 108.055 31.935 108.875 ;
        RECT 32.145 108.730 32.315 109.530 ;
        RECT 32.600 109.505 33.265 109.675 ;
        RECT 34.445 109.530 34.715 110.435 ;
        RECT 34.885 109.845 35.215 110.605 ;
        RECT 35.395 109.675 35.565 110.435 ;
        RECT 32.600 109.360 32.770 109.505 ;
        RECT 32.485 109.030 32.770 109.360 ;
        RECT 32.600 108.775 32.770 109.030 ;
        RECT 33.005 108.955 33.335 109.325 ;
        RECT 32.145 108.225 32.405 108.730 ;
        RECT 32.600 108.605 33.265 108.775 ;
        RECT 32.585 108.055 32.915 108.435 ;
        RECT 33.095 108.225 33.265 108.605 ;
        RECT 34.445 108.730 34.615 109.530 ;
        RECT 34.900 109.505 35.565 109.675 ;
        RECT 36.285 109.515 38.875 110.605 ;
        RECT 39.050 110.170 44.395 110.605 ;
        RECT 44.570 110.170 49.915 110.605 ;
        RECT 34.900 109.360 35.070 109.505 ;
        RECT 34.785 109.030 35.070 109.360 ;
        RECT 34.900 108.775 35.070 109.030 ;
        RECT 35.305 108.955 35.635 109.325 ;
        RECT 36.285 108.995 37.495 109.515 ;
        RECT 37.665 108.825 38.875 109.345 ;
        RECT 40.640 108.920 40.990 110.170 ;
        RECT 34.445 108.225 34.705 108.730 ;
        RECT 34.900 108.605 35.565 108.775 ;
        RECT 34.885 108.055 35.215 108.435 ;
        RECT 35.395 108.225 35.565 108.605 ;
        RECT 36.285 108.055 38.875 108.825 ;
        RECT 42.470 108.600 42.810 109.430 ;
        RECT 46.160 108.920 46.510 110.170 ;
        RECT 50.085 109.440 50.375 110.605 ;
        RECT 51.095 109.675 51.265 110.435 ;
        RECT 51.445 109.845 51.775 110.605 ;
        RECT 51.095 109.505 51.760 109.675 ;
        RECT 51.945 109.530 52.215 110.435 ;
        RECT 47.990 108.600 48.330 109.430 ;
        RECT 51.590 109.360 51.760 109.505 ;
        RECT 51.025 108.955 51.355 109.325 ;
        RECT 51.590 109.030 51.875 109.360 ;
        RECT 39.050 108.055 44.395 108.600 ;
        RECT 44.570 108.055 49.915 108.600 ;
        RECT 50.085 108.055 50.375 108.780 ;
        RECT 51.590 108.775 51.760 109.030 ;
        RECT 51.095 108.605 51.760 108.775 ;
        RECT 52.045 108.730 52.215 109.530 ;
        RECT 53.305 109.515 56.815 110.605 ;
        RECT 57.075 109.675 57.245 110.435 ;
        RECT 57.425 109.845 57.755 110.605 ;
        RECT 53.305 108.995 54.995 109.515 ;
        RECT 57.075 109.505 57.740 109.675 ;
        RECT 57.925 109.530 58.195 110.435 ;
        RECT 57.570 109.360 57.740 109.505 ;
        RECT 55.165 108.825 56.815 109.345 ;
        RECT 57.005 108.955 57.335 109.325 ;
        RECT 57.570 109.030 57.855 109.360 ;
        RECT 51.095 108.225 51.265 108.605 ;
        RECT 51.445 108.055 51.775 108.435 ;
        RECT 51.955 108.225 52.215 108.730 ;
        RECT 53.305 108.055 56.815 108.825 ;
        RECT 57.570 108.775 57.740 109.030 ;
        RECT 57.075 108.605 57.740 108.775 ;
        RECT 58.025 108.730 58.195 109.530 ;
        RECT 58.365 109.515 59.575 110.605 ;
        RECT 59.755 109.625 60.085 110.435 ;
        RECT 60.255 109.805 60.495 110.605 ;
        RECT 58.365 108.975 58.885 109.515 ;
        RECT 59.755 109.455 60.470 109.625 ;
        RECT 59.055 108.805 59.575 109.345 ;
        RECT 59.750 109.045 60.130 109.285 ;
        RECT 60.300 109.215 60.470 109.455 ;
        RECT 60.675 109.585 60.845 110.435 ;
        RECT 61.015 109.805 61.345 110.605 ;
        RECT 61.515 109.585 61.685 110.435 ;
        RECT 60.675 109.415 61.685 109.585 ;
        RECT 61.855 109.455 62.185 110.605 ;
        RECT 62.965 109.515 64.635 110.605 ;
        RECT 61.190 109.245 61.685 109.415 ;
        RECT 60.300 109.045 60.800 109.215 ;
        RECT 61.185 109.075 61.685 109.245 ;
        RECT 60.300 108.875 60.470 109.045 ;
        RECT 61.190 108.875 61.685 109.075 ;
        RECT 62.965 108.995 63.715 109.515 ;
        RECT 64.845 109.465 65.075 110.605 ;
        RECT 65.245 109.455 65.575 110.435 ;
        RECT 65.745 109.465 65.955 110.605 ;
        RECT 66.645 109.515 68.315 110.605 ;
        RECT 68.575 109.675 68.745 110.435 ;
        RECT 68.925 109.845 69.255 110.605 ;
        RECT 57.075 108.225 57.245 108.605 ;
        RECT 57.425 108.055 57.755 108.435 ;
        RECT 57.935 108.225 58.195 108.730 ;
        RECT 58.365 108.055 59.575 108.805 ;
        RECT 59.835 108.705 60.470 108.875 ;
        RECT 60.675 108.705 61.685 108.875 ;
        RECT 59.835 108.225 60.005 108.705 ;
        RECT 60.185 108.055 60.425 108.535 ;
        RECT 60.675 108.225 60.845 108.705 ;
        RECT 61.015 108.055 61.345 108.535 ;
        RECT 61.515 108.225 61.685 108.705 ;
        RECT 61.855 108.055 62.185 108.855 ;
        RECT 63.885 108.825 64.635 109.345 ;
        RECT 64.825 109.045 65.155 109.295 ;
        RECT 62.965 108.055 64.635 108.825 ;
        RECT 64.845 108.055 65.075 108.875 ;
        RECT 65.325 108.855 65.575 109.455 ;
        RECT 66.645 108.995 67.395 109.515 ;
        RECT 68.575 109.505 69.240 109.675 ;
        RECT 69.425 109.530 69.695 110.435 ;
        RECT 70.330 110.170 75.675 110.605 ;
        RECT 69.070 109.360 69.240 109.505 ;
        RECT 65.245 108.225 65.575 108.855 ;
        RECT 65.745 108.055 65.955 108.875 ;
        RECT 67.565 108.825 68.315 109.345 ;
        RECT 68.505 108.955 68.835 109.325 ;
        RECT 69.070 109.030 69.355 109.360 ;
        RECT 66.645 108.055 68.315 108.825 ;
        RECT 69.070 108.775 69.240 109.030 ;
        RECT 68.575 108.605 69.240 108.775 ;
        RECT 69.525 108.730 69.695 109.530 ;
        RECT 71.920 108.920 72.270 110.170 ;
        RECT 75.845 109.440 76.135 110.605 ;
        RECT 76.365 109.465 76.575 110.605 ;
        RECT 76.745 109.455 77.075 110.435 ;
        RECT 77.245 109.465 77.475 110.605 ;
        RECT 77.745 109.465 77.955 110.605 ;
        RECT 78.125 109.455 78.455 110.435 ;
        RECT 78.625 109.465 78.855 110.605 ;
        RECT 79.995 109.625 80.325 110.435 ;
        RECT 80.495 109.805 80.735 110.605 ;
        RECT 79.995 109.455 80.710 109.625 ;
        RECT 68.575 108.225 68.745 108.605 ;
        RECT 68.925 108.055 69.255 108.435 ;
        RECT 69.435 108.225 69.695 108.730 ;
        RECT 73.750 108.600 74.090 109.430 ;
        RECT 70.330 108.055 75.675 108.600 ;
        RECT 75.845 108.055 76.135 108.780 ;
        RECT 76.365 108.055 76.575 108.875 ;
        RECT 76.745 108.855 76.995 109.455 ;
        RECT 77.165 109.045 77.495 109.295 ;
        RECT 76.745 108.225 77.075 108.855 ;
        RECT 77.245 108.055 77.475 108.875 ;
        RECT 77.745 108.055 77.955 108.875 ;
        RECT 78.125 108.855 78.375 109.455 ;
        RECT 78.545 109.045 78.875 109.295 ;
        RECT 79.990 109.045 80.370 109.285 ;
        RECT 80.540 109.215 80.710 109.455 ;
        RECT 80.915 109.585 81.085 110.435 ;
        RECT 81.255 109.805 81.585 110.605 ;
        RECT 81.755 109.585 81.925 110.435 ;
        RECT 80.915 109.415 81.925 109.585 ;
        RECT 82.095 109.455 82.425 110.605 ;
        RECT 82.835 109.675 83.005 110.435 ;
        RECT 83.185 109.845 83.515 110.605 ;
        RECT 82.835 109.505 83.500 109.675 ;
        RECT 83.685 109.530 83.955 110.435 ;
        RECT 80.540 109.045 81.040 109.215 ;
        RECT 80.540 108.875 80.710 109.045 ;
        RECT 81.430 108.875 81.925 109.415 ;
        RECT 83.330 109.360 83.500 109.505 ;
        RECT 82.765 108.955 83.095 109.325 ;
        RECT 83.330 109.030 83.615 109.360 ;
        RECT 78.125 108.225 78.455 108.855 ;
        RECT 78.625 108.055 78.855 108.875 ;
        RECT 80.075 108.705 80.710 108.875 ;
        RECT 80.915 108.705 81.925 108.875 ;
        RECT 80.075 108.225 80.245 108.705 ;
        RECT 80.425 108.055 80.665 108.535 ;
        RECT 80.915 108.225 81.085 108.705 ;
        RECT 81.255 108.055 81.585 108.535 ;
        RECT 81.755 108.225 81.925 108.705 ;
        RECT 82.095 108.055 82.425 108.855 ;
        RECT 83.330 108.775 83.500 109.030 ;
        RECT 82.835 108.605 83.500 108.775 ;
        RECT 83.785 108.730 83.955 109.530 ;
        RECT 84.585 109.515 87.175 110.605 ;
        RECT 84.585 108.995 85.795 109.515 ;
        RECT 87.385 109.465 87.615 110.605 ;
        RECT 87.785 109.455 88.115 110.435 ;
        RECT 88.285 109.465 88.495 110.605 ;
        RECT 88.725 109.515 92.235 110.605 ;
        RECT 85.965 108.825 87.175 109.345 ;
        RECT 87.365 109.045 87.695 109.295 ;
        RECT 82.835 108.225 83.005 108.605 ;
        RECT 83.185 108.055 83.515 108.435 ;
        RECT 83.695 108.225 83.955 108.730 ;
        RECT 84.585 108.055 87.175 108.825 ;
        RECT 87.385 108.055 87.615 108.875 ;
        RECT 87.865 108.855 88.115 109.455 ;
        RECT 88.725 108.995 90.415 109.515 ;
        RECT 92.445 109.465 92.675 110.605 ;
        RECT 92.845 109.455 93.175 110.435 ;
        RECT 93.345 109.465 93.555 110.605 ;
        RECT 93.875 109.675 94.045 110.435 ;
        RECT 94.225 109.845 94.555 110.605 ;
        RECT 93.875 109.505 94.540 109.675 ;
        RECT 94.725 109.530 94.995 110.435 ;
        RECT 87.785 108.225 88.115 108.855 ;
        RECT 88.285 108.055 88.495 108.875 ;
        RECT 90.585 108.825 92.235 109.345 ;
        RECT 92.425 109.045 92.755 109.295 ;
        RECT 88.725 108.055 92.235 108.825 ;
        RECT 92.445 108.055 92.675 108.875 ;
        RECT 92.925 108.855 93.175 109.455 ;
        RECT 94.370 109.360 94.540 109.505 ;
        RECT 93.805 108.955 94.135 109.325 ;
        RECT 94.370 109.030 94.655 109.360 ;
        RECT 92.845 108.225 93.175 108.855 ;
        RECT 93.345 108.055 93.555 108.875 ;
        RECT 94.370 108.775 94.540 109.030 ;
        RECT 93.875 108.605 94.540 108.775 ;
        RECT 94.825 108.730 94.995 109.530 ;
        RECT 95.165 109.515 96.375 110.605 ;
        RECT 96.545 109.515 100.055 110.605 ;
        RECT 100.225 109.530 100.495 110.435 ;
        RECT 100.665 109.845 100.995 110.605 ;
        RECT 101.175 109.675 101.345 110.435 ;
        RECT 95.165 108.975 95.685 109.515 ;
        RECT 95.855 108.805 96.375 109.345 ;
        RECT 96.545 108.995 98.235 109.515 ;
        RECT 98.405 108.825 100.055 109.345 ;
        RECT 93.875 108.225 94.045 108.605 ;
        RECT 94.225 108.055 94.555 108.435 ;
        RECT 94.735 108.225 94.995 108.730 ;
        RECT 95.165 108.055 96.375 108.805 ;
        RECT 96.545 108.055 100.055 108.825 ;
        RECT 100.225 108.730 100.395 109.530 ;
        RECT 100.680 109.505 101.345 109.675 ;
        RECT 100.680 109.360 100.850 109.505 ;
        RECT 101.605 109.440 101.895 110.605 ;
        RECT 102.525 109.515 106.035 110.605 ;
        RECT 106.295 109.675 106.465 110.435 ;
        RECT 106.645 109.845 106.975 110.605 ;
        RECT 100.565 109.030 100.850 109.360 ;
        RECT 100.680 108.775 100.850 109.030 ;
        RECT 101.085 108.955 101.415 109.325 ;
        RECT 102.525 108.995 104.215 109.515 ;
        RECT 106.295 109.505 106.960 109.675 ;
        RECT 107.145 109.530 107.415 110.435 ;
        RECT 106.790 109.360 106.960 109.505 ;
        RECT 104.385 108.825 106.035 109.345 ;
        RECT 106.225 108.955 106.555 109.325 ;
        RECT 106.790 109.030 107.075 109.360 ;
        RECT 100.225 108.225 100.485 108.730 ;
        RECT 100.680 108.605 101.345 108.775 ;
        RECT 100.665 108.055 100.995 108.435 ;
        RECT 101.175 108.225 101.345 108.605 ;
        RECT 101.605 108.055 101.895 108.780 ;
        RECT 102.525 108.055 106.035 108.825 ;
        RECT 106.790 108.775 106.960 109.030 ;
        RECT 106.295 108.605 106.960 108.775 ;
        RECT 107.245 108.730 107.415 109.530 ;
        RECT 107.585 109.515 108.795 110.605 ;
        RECT 107.585 108.975 108.105 109.515 ;
        RECT 109.025 109.465 109.235 110.605 ;
        RECT 109.405 109.455 109.735 110.435 ;
        RECT 109.905 109.465 110.135 110.605 ;
        RECT 110.435 109.675 110.605 110.435 ;
        RECT 110.785 109.845 111.115 110.605 ;
        RECT 110.435 109.505 111.100 109.675 ;
        RECT 111.285 109.530 111.555 110.435 ;
        RECT 108.275 108.805 108.795 109.345 ;
        RECT 106.295 108.225 106.465 108.605 ;
        RECT 106.645 108.055 106.975 108.435 ;
        RECT 107.155 108.225 107.415 108.730 ;
        RECT 107.585 108.055 108.795 108.805 ;
        RECT 109.025 108.055 109.235 108.875 ;
        RECT 109.405 108.855 109.655 109.455 ;
        RECT 110.930 109.360 111.100 109.505 ;
        RECT 109.825 109.045 110.155 109.295 ;
        RECT 110.365 108.955 110.695 109.325 ;
        RECT 110.930 109.030 111.215 109.360 ;
        RECT 109.405 108.225 109.735 108.855 ;
        RECT 109.905 108.055 110.135 108.875 ;
        RECT 110.930 108.775 111.100 109.030 ;
        RECT 110.435 108.605 111.100 108.775 ;
        RECT 111.385 108.730 111.555 109.530 ;
        RECT 111.815 109.675 111.985 110.435 ;
        RECT 112.165 109.845 112.495 110.605 ;
        RECT 111.815 109.505 112.480 109.675 ;
        RECT 112.665 109.530 112.935 110.435 ;
        RECT 112.310 109.360 112.480 109.505 ;
        RECT 111.745 108.955 112.075 109.325 ;
        RECT 112.310 109.030 112.595 109.360 ;
        RECT 112.310 108.775 112.480 109.030 ;
        RECT 110.435 108.225 110.605 108.605 ;
        RECT 110.785 108.055 111.115 108.435 ;
        RECT 111.295 108.225 111.555 108.730 ;
        RECT 111.815 108.605 112.480 108.775 ;
        RECT 112.765 108.730 112.935 109.530 ;
        RECT 113.105 109.515 114.315 110.605 ;
        RECT 113.105 108.975 113.625 109.515 ;
        RECT 114.525 109.465 114.755 110.605 ;
        RECT 114.925 109.455 115.255 110.435 ;
        RECT 115.425 109.465 115.635 110.605 ;
        RECT 115.870 109.935 116.125 110.435 ;
        RECT 116.295 110.105 116.625 110.605 ;
        RECT 115.870 109.765 116.620 109.935 ;
        RECT 113.795 108.805 114.315 109.345 ;
        RECT 114.505 109.045 114.835 109.295 ;
        RECT 111.815 108.225 111.985 108.605 ;
        RECT 112.165 108.055 112.495 108.435 ;
        RECT 112.675 108.225 112.935 108.730 ;
        RECT 113.105 108.055 114.315 108.805 ;
        RECT 114.525 108.055 114.755 108.875 ;
        RECT 115.005 108.855 115.255 109.455 ;
        RECT 115.870 108.945 116.220 109.595 ;
        RECT 114.925 108.225 115.255 108.855 ;
        RECT 115.425 108.055 115.635 108.875 ;
        RECT 116.390 108.775 116.620 109.765 ;
        RECT 115.870 108.605 116.620 108.775 ;
        RECT 115.870 108.315 116.125 108.605 ;
        RECT 116.295 108.055 116.625 108.435 ;
        RECT 116.795 108.315 116.965 110.435 ;
        RECT 117.135 109.635 117.460 110.420 ;
        RECT 117.630 110.145 117.880 110.605 ;
        RECT 118.050 110.105 118.300 110.435 ;
        RECT 118.515 110.105 119.195 110.435 ;
        RECT 118.050 109.975 118.220 110.105 ;
        RECT 117.825 109.805 118.220 109.975 ;
        RECT 117.195 108.585 117.655 109.635 ;
        RECT 117.825 108.445 117.995 109.805 ;
        RECT 118.390 109.545 118.855 109.935 ;
        RECT 118.165 108.735 118.515 109.355 ;
        RECT 118.685 108.955 118.855 109.545 ;
        RECT 119.025 109.325 119.195 110.105 ;
        RECT 119.365 110.005 119.535 110.345 ;
        RECT 119.770 110.175 120.100 110.605 ;
        RECT 120.270 110.005 120.440 110.345 ;
        RECT 120.735 110.145 121.105 110.605 ;
        RECT 119.365 109.835 120.440 110.005 ;
        RECT 121.275 109.975 121.445 110.435 ;
        RECT 121.680 110.095 122.550 110.435 ;
        RECT 122.720 110.145 122.970 110.605 ;
        RECT 120.885 109.805 121.445 109.975 ;
        RECT 120.885 109.665 121.055 109.805 ;
        RECT 119.555 109.495 121.055 109.665 ;
        RECT 121.750 109.635 122.210 109.925 ;
        RECT 119.025 109.155 120.715 109.325 ;
        RECT 118.685 108.735 119.040 108.955 ;
        RECT 119.210 108.445 119.380 109.155 ;
        RECT 119.585 108.735 120.375 108.985 ;
        RECT 120.545 108.975 120.715 109.155 ;
        RECT 120.885 108.805 121.055 109.495 ;
        RECT 117.325 108.055 117.655 108.415 ;
        RECT 117.825 108.275 118.320 108.445 ;
        RECT 118.525 108.275 119.380 108.445 ;
        RECT 120.255 108.055 120.585 108.515 ;
        RECT 120.795 108.415 121.055 108.805 ;
        RECT 121.245 109.625 122.210 109.635 ;
        RECT 122.380 109.715 122.550 110.095 ;
        RECT 123.140 110.055 123.310 110.345 ;
        RECT 123.490 110.225 123.820 110.605 ;
        RECT 123.140 109.885 123.940 110.055 ;
        RECT 121.245 109.465 121.920 109.625 ;
        RECT 122.380 109.545 123.600 109.715 ;
        RECT 121.245 108.675 121.455 109.465 ;
        RECT 122.380 109.455 122.550 109.545 ;
        RECT 121.625 108.675 121.975 109.295 ;
        RECT 122.145 109.285 122.550 109.455 ;
        RECT 122.145 108.505 122.315 109.285 ;
        RECT 122.485 108.835 122.705 109.115 ;
        RECT 122.885 109.005 123.425 109.375 ;
        RECT 123.770 109.265 123.940 109.885 ;
        RECT 124.115 109.545 124.285 110.605 ;
        RECT 124.495 109.595 124.785 110.435 ;
        RECT 124.955 109.765 125.125 110.605 ;
        RECT 125.335 109.595 125.585 110.435 ;
        RECT 125.795 109.765 125.965 110.605 ;
        RECT 124.495 109.425 126.220 109.595 ;
        RECT 122.485 108.665 123.015 108.835 ;
        RECT 120.795 108.245 121.145 108.415 ;
        RECT 121.365 108.225 122.315 108.505 ;
        RECT 122.485 108.055 122.675 108.495 ;
        RECT 122.845 108.435 123.015 108.665 ;
        RECT 123.185 108.605 123.425 109.005 ;
        RECT 123.595 109.255 123.940 109.265 ;
        RECT 123.595 109.045 125.625 109.255 ;
        RECT 123.595 108.790 123.920 109.045 ;
        RECT 125.810 108.875 126.220 109.425 ;
        RECT 126.445 109.515 127.655 110.605 ;
        RECT 126.445 108.975 126.965 109.515 ;
        RECT 123.595 108.435 123.915 108.790 ;
        RECT 122.845 108.265 123.915 108.435 ;
        RECT 124.115 108.055 124.285 108.865 ;
        RECT 124.455 108.705 126.220 108.875 ;
        RECT 127.135 108.805 127.655 109.345 ;
        RECT 124.455 108.225 124.785 108.705 ;
        RECT 124.955 108.055 125.125 108.525 ;
        RECT 125.295 108.225 125.625 108.705 ;
        RECT 125.795 108.055 125.965 108.525 ;
        RECT 126.445 108.055 127.655 108.805 ;
        RECT 14.580 107.885 127.740 108.055 ;
        RECT 14.665 107.135 15.875 107.885 ;
        RECT 16.355 107.415 16.525 107.885 ;
        RECT 16.695 107.235 17.025 107.715 ;
        RECT 17.195 107.415 17.365 107.885 ;
        RECT 17.535 107.235 17.865 107.715 ;
        RECT 14.665 106.595 15.185 107.135 ;
        RECT 16.100 107.065 17.865 107.235 ;
        RECT 18.035 107.075 18.205 107.885 ;
        RECT 18.405 107.505 19.475 107.675 ;
        RECT 18.405 107.150 18.725 107.505 ;
        RECT 15.355 106.425 15.875 106.965 ;
        RECT 14.665 105.335 15.875 106.425 ;
        RECT 16.100 106.515 16.510 107.065 ;
        RECT 18.400 106.895 18.725 107.150 ;
        RECT 16.695 106.685 18.725 106.895 ;
        RECT 18.380 106.675 18.725 106.685 ;
        RECT 18.895 106.935 19.135 107.335 ;
        RECT 19.305 107.275 19.475 107.505 ;
        RECT 19.645 107.445 19.835 107.885 ;
        RECT 20.005 107.435 20.955 107.715 ;
        RECT 21.175 107.525 21.525 107.695 ;
        RECT 19.305 107.105 19.835 107.275 ;
        RECT 16.100 106.345 17.825 106.515 ;
        RECT 16.355 105.335 16.525 106.175 ;
        RECT 16.735 105.505 16.985 106.345 ;
        RECT 17.195 105.335 17.365 106.175 ;
        RECT 17.535 105.505 17.825 106.345 ;
        RECT 18.035 105.335 18.205 106.395 ;
        RECT 18.380 106.055 18.550 106.675 ;
        RECT 18.895 106.565 19.435 106.935 ;
        RECT 19.615 106.825 19.835 107.105 ;
        RECT 20.005 106.655 20.175 107.435 ;
        RECT 19.770 106.485 20.175 106.655 ;
        RECT 20.345 106.645 20.695 107.265 ;
        RECT 19.770 106.395 19.940 106.485 ;
        RECT 20.865 106.475 21.075 107.265 ;
        RECT 18.720 106.225 19.940 106.395 ;
        RECT 20.400 106.315 21.075 106.475 ;
        RECT 18.380 105.885 19.180 106.055 ;
        RECT 18.500 105.335 18.830 105.715 ;
        RECT 19.010 105.595 19.180 105.885 ;
        RECT 19.770 105.845 19.940 106.225 ;
        RECT 20.110 106.305 21.075 106.315 ;
        RECT 21.265 107.135 21.525 107.525 ;
        RECT 21.735 107.425 22.065 107.885 ;
        RECT 22.940 107.495 23.795 107.665 ;
        RECT 24.000 107.495 24.495 107.665 ;
        RECT 24.665 107.525 24.995 107.885 ;
        RECT 21.265 106.445 21.435 107.135 ;
        RECT 21.605 106.785 21.775 106.965 ;
        RECT 21.945 106.955 22.735 107.205 ;
        RECT 22.940 106.785 23.110 107.495 ;
        RECT 23.280 106.985 23.635 107.205 ;
        RECT 21.605 106.615 23.295 106.785 ;
        RECT 20.110 106.015 20.570 106.305 ;
        RECT 21.265 106.275 22.765 106.445 ;
        RECT 21.265 106.135 21.435 106.275 ;
        RECT 20.875 105.965 21.435 106.135 ;
        RECT 19.350 105.335 19.600 105.795 ;
        RECT 19.770 105.505 20.640 105.845 ;
        RECT 20.875 105.505 21.045 105.965 ;
        RECT 21.880 105.935 22.955 106.105 ;
        RECT 21.215 105.335 21.585 105.795 ;
        RECT 21.880 105.595 22.050 105.935 ;
        RECT 22.220 105.335 22.550 105.765 ;
        RECT 22.785 105.595 22.955 105.935 ;
        RECT 23.125 105.835 23.295 106.615 ;
        RECT 23.465 106.395 23.635 106.985 ;
        RECT 23.805 106.585 24.155 107.205 ;
        RECT 23.465 106.005 23.930 106.395 ;
        RECT 24.325 106.135 24.495 107.495 ;
        RECT 24.665 106.305 25.125 107.355 ;
        RECT 24.100 105.965 24.495 106.135 ;
        RECT 24.100 105.835 24.270 105.965 ;
        RECT 23.125 105.505 23.805 105.835 ;
        RECT 24.020 105.505 24.270 105.835 ;
        RECT 24.440 105.335 24.690 105.795 ;
        RECT 24.860 105.520 25.185 106.305 ;
        RECT 25.355 105.505 25.525 107.625 ;
        RECT 25.695 107.505 26.025 107.885 ;
        RECT 26.195 107.335 26.450 107.625 ;
        RECT 26.935 107.415 27.105 107.885 ;
        RECT 25.700 107.165 26.450 107.335 ;
        RECT 27.275 107.235 27.605 107.715 ;
        RECT 27.775 107.415 27.945 107.885 ;
        RECT 28.115 107.235 28.445 107.715 ;
        RECT 25.700 106.175 25.930 107.165 ;
        RECT 26.680 107.065 28.445 107.235 ;
        RECT 28.615 107.075 28.785 107.885 ;
        RECT 28.985 107.505 30.055 107.675 ;
        RECT 28.985 107.150 29.305 107.505 ;
        RECT 26.100 106.345 26.450 106.995 ;
        RECT 26.680 106.515 27.090 107.065 ;
        RECT 28.980 106.895 29.305 107.150 ;
        RECT 27.275 106.685 29.305 106.895 ;
        RECT 28.960 106.675 29.305 106.685 ;
        RECT 29.475 106.935 29.715 107.335 ;
        RECT 29.885 107.275 30.055 107.505 ;
        RECT 30.225 107.445 30.415 107.885 ;
        RECT 30.585 107.435 31.535 107.715 ;
        RECT 31.755 107.525 32.105 107.695 ;
        RECT 29.885 107.105 30.415 107.275 ;
        RECT 26.680 106.345 28.405 106.515 ;
        RECT 25.700 106.005 26.450 106.175 ;
        RECT 25.695 105.335 26.025 105.835 ;
        RECT 26.195 105.505 26.450 106.005 ;
        RECT 26.935 105.335 27.105 106.175 ;
        RECT 27.315 105.505 27.565 106.345 ;
        RECT 27.775 105.335 27.945 106.175 ;
        RECT 28.115 105.505 28.405 106.345 ;
        RECT 28.615 105.335 28.785 106.395 ;
        RECT 28.960 106.055 29.130 106.675 ;
        RECT 29.475 106.565 30.015 106.935 ;
        RECT 30.195 106.825 30.415 107.105 ;
        RECT 30.585 106.655 30.755 107.435 ;
        RECT 30.350 106.485 30.755 106.655 ;
        RECT 30.925 106.645 31.275 107.265 ;
        RECT 30.350 106.395 30.520 106.485 ;
        RECT 31.445 106.475 31.655 107.265 ;
        RECT 29.300 106.225 30.520 106.395 ;
        RECT 30.980 106.315 31.655 106.475 ;
        RECT 28.960 105.885 29.760 106.055 ;
        RECT 29.080 105.335 29.410 105.715 ;
        RECT 29.590 105.595 29.760 105.885 ;
        RECT 30.350 105.845 30.520 106.225 ;
        RECT 30.690 106.305 31.655 106.315 ;
        RECT 31.845 107.135 32.105 107.525 ;
        RECT 32.315 107.425 32.645 107.885 ;
        RECT 33.520 107.495 34.375 107.665 ;
        RECT 34.580 107.495 35.075 107.665 ;
        RECT 35.245 107.525 35.575 107.885 ;
        RECT 31.845 106.445 32.015 107.135 ;
        RECT 32.185 106.785 32.355 106.965 ;
        RECT 32.525 106.955 33.315 107.205 ;
        RECT 33.520 106.785 33.690 107.495 ;
        RECT 33.860 106.985 34.215 107.205 ;
        RECT 32.185 106.615 33.875 106.785 ;
        RECT 30.690 106.015 31.150 106.305 ;
        RECT 31.845 106.275 33.345 106.445 ;
        RECT 31.845 106.135 32.015 106.275 ;
        RECT 31.455 105.965 32.015 106.135 ;
        RECT 29.930 105.335 30.180 105.795 ;
        RECT 30.350 105.505 31.220 105.845 ;
        RECT 31.455 105.505 31.625 105.965 ;
        RECT 32.460 105.935 33.535 106.105 ;
        RECT 31.795 105.335 32.165 105.795 ;
        RECT 32.460 105.595 32.630 105.935 ;
        RECT 32.800 105.335 33.130 105.765 ;
        RECT 33.365 105.595 33.535 105.935 ;
        RECT 33.705 105.835 33.875 106.615 ;
        RECT 34.045 106.395 34.215 106.985 ;
        RECT 34.385 106.585 34.735 107.205 ;
        RECT 34.045 106.005 34.510 106.395 ;
        RECT 34.905 106.135 35.075 107.495 ;
        RECT 35.245 106.305 35.705 107.355 ;
        RECT 34.680 105.965 35.075 106.135 ;
        RECT 34.680 105.835 34.850 105.965 ;
        RECT 33.705 105.505 34.385 105.835 ;
        RECT 34.600 105.505 34.850 105.835 ;
        RECT 35.020 105.335 35.270 105.795 ;
        RECT 35.440 105.520 35.765 106.305 ;
        RECT 35.935 105.505 36.105 107.625 ;
        RECT 36.275 107.505 36.605 107.885 ;
        RECT 36.775 107.335 37.030 107.625 ;
        RECT 36.280 107.165 37.030 107.335 ;
        RECT 36.280 106.175 36.510 107.165 ;
        RECT 37.205 107.160 37.495 107.885 ;
        RECT 37.665 107.210 37.925 107.715 ;
        RECT 38.105 107.505 38.435 107.885 ;
        RECT 38.615 107.335 38.785 107.715 ;
        RECT 36.680 106.345 37.030 106.995 ;
        RECT 36.280 106.005 37.030 106.175 ;
        RECT 36.275 105.335 36.605 105.835 ;
        RECT 36.775 105.505 37.030 106.005 ;
        RECT 37.205 105.335 37.495 106.500 ;
        RECT 37.665 106.410 37.835 107.210 ;
        RECT 38.120 107.165 38.785 107.335 ;
        RECT 38.120 106.910 38.290 107.165 ;
        RECT 39.565 107.065 39.775 107.885 ;
        RECT 39.945 107.085 40.275 107.715 ;
        RECT 38.005 106.580 38.290 106.910 ;
        RECT 38.525 106.615 38.855 106.985 ;
        RECT 38.120 106.435 38.290 106.580 ;
        RECT 39.945 106.485 40.195 107.085 ;
        RECT 40.445 107.065 40.675 107.885 ;
        RECT 40.885 107.135 42.095 107.885 ;
        RECT 40.365 106.645 40.695 106.895 ;
        RECT 37.665 105.505 37.935 106.410 ;
        RECT 38.120 106.265 38.785 106.435 ;
        RECT 38.105 105.335 38.435 106.095 ;
        RECT 38.615 105.505 38.785 106.265 ;
        RECT 39.565 105.335 39.775 106.475 ;
        RECT 39.945 105.505 40.275 106.485 ;
        RECT 40.445 105.335 40.675 106.475 ;
        RECT 40.885 106.425 41.405 106.965 ;
        RECT 41.575 106.595 42.095 107.135 ;
        RECT 42.265 107.210 42.525 107.715 ;
        RECT 42.705 107.505 43.035 107.885 ;
        RECT 43.215 107.335 43.385 107.715 ;
        RECT 40.885 105.335 42.095 106.425 ;
        RECT 42.265 106.410 42.435 107.210 ;
        RECT 42.720 107.165 43.385 107.335 ;
        RECT 42.720 106.910 42.890 107.165 ;
        RECT 44.165 107.065 44.375 107.885 ;
        RECT 44.545 107.085 44.875 107.715 ;
        RECT 42.605 106.580 42.890 106.910 ;
        RECT 43.125 106.615 43.455 106.985 ;
        RECT 42.720 106.435 42.890 106.580 ;
        RECT 44.545 106.485 44.795 107.085 ;
        RECT 45.045 107.065 45.275 107.885 ;
        RECT 45.575 107.335 45.745 107.715 ;
        RECT 45.925 107.505 46.255 107.885 ;
        RECT 45.575 107.165 46.240 107.335 ;
        RECT 46.435 107.210 46.695 107.715 ;
        RECT 47.175 107.415 47.345 107.885 ;
        RECT 47.515 107.235 47.845 107.715 ;
        RECT 48.015 107.415 48.185 107.885 ;
        RECT 48.355 107.235 48.685 107.715 ;
        RECT 44.965 106.645 45.295 106.895 ;
        RECT 45.505 106.615 45.835 106.985 ;
        RECT 46.070 106.910 46.240 107.165 ;
        RECT 46.070 106.580 46.355 106.910 ;
        RECT 42.265 105.505 42.535 106.410 ;
        RECT 42.720 106.265 43.385 106.435 ;
        RECT 42.705 105.335 43.035 106.095 ;
        RECT 43.215 105.505 43.385 106.265 ;
        RECT 44.165 105.335 44.375 106.475 ;
        RECT 44.545 105.505 44.875 106.485 ;
        RECT 45.045 105.335 45.275 106.475 ;
        RECT 46.070 106.435 46.240 106.580 ;
        RECT 45.575 106.265 46.240 106.435 ;
        RECT 46.525 106.410 46.695 107.210 ;
        RECT 45.575 105.505 45.745 106.265 ;
        RECT 45.925 105.335 46.255 106.095 ;
        RECT 46.425 105.505 46.695 106.410 ;
        RECT 46.920 107.065 48.685 107.235 ;
        RECT 48.855 107.075 49.025 107.885 ;
        RECT 49.225 107.505 50.295 107.675 ;
        RECT 49.225 107.150 49.545 107.505 ;
        RECT 46.920 106.515 47.330 107.065 ;
        RECT 49.220 106.895 49.545 107.150 ;
        RECT 47.515 106.685 49.545 106.895 ;
        RECT 49.200 106.675 49.545 106.685 ;
        RECT 49.715 106.935 49.955 107.335 ;
        RECT 50.125 107.275 50.295 107.505 ;
        RECT 50.465 107.445 50.655 107.885 ;
        RECT 50.825 107.435 51.775 107.715 ;
        RECT 51.995 107.525 52.345 107.695 ;
        RECT 50.125 107.105 50.655 107.275 ;
        RECT 46.920 106.345 48.645 106.515 ;
        RECT 47.175 105.335 47.345 106.175 ;
        RECT 47.555 105.505 47.805 106.345 ;
        RECT 48.015 105.335 48.185 106.175 ;
        RECT 48.355 105.505 48.645 106.345 ;
        RECT 48.855 105.335 49.025 106.395 ;
        RECT 49.200 106.055 49.370 106.675 ;
        RECT 49.715 106.565 50.255 106.935 ;
        RECT 50.435 106.825 50.655 107.105 ;
        RECT 50.825 106.655 50.995 107.435 ;
        RECT 50.590 106.485 50.995 106.655 ;
        RECT 51.165 106.645 51.515 107.265 ;
        RECT 50.590 106.395 50.760 106.485 ;
        RECT 51.685 106.475 51.895 107.265 ;
        RECT 49.540 106.225 50.760 106.395 ;
        RECT 51.220 106.315 51.895 106.475 ;
        RECT 49.200 105.885 50.000 106.055 ;
        RECT 49.320 105.335 49.650 105.715 ;
        RECT 49.830 105.595 50.000 105.885 ;
        RECT 50.590 105.845 50.760 106.225 ;
        RECT 50.930 106.305 51.895 106.315 ;
        RECT 52.085 107.135 52.345 107.525 ;
        RECT 52.555 107.425 52.885 107.885 ;
        RECT 53.760 107.495 54.615 107.665 ;
        RECT 54.820 107.495 55.315 107.665 ;
        RECT 55.485 107.525 55.815 107.885 ;
        RECT 52.085 106.445 52.255 107.135 ;
        RECT 52.425 106.785 52.595 106.965 ;
        RECT 52.765 106.955 53.555 107.205 ;
        RECT 53.760 106.785 53.930 107.495 ;
        RECT 54.100 106.985 54.455 107.205 ;
        RECT 52.425 106.615 54.115 106.785 ;
        RECT 50.930 106.015 51.390 106.305 ;
        RECT 52.085 106.275 53.585 106.445 ;
        RECT 52.085 106.135 52.255 106.275 ;
        RECT 51.695 105.965 52.255 106.135 ;
        RECT 50.170 105.335 50.420 105.795 ;
        RECT 50.590 105.505 51.460 105.845 ;
        RECT 51.695 105.505 51.865 105.965 ;
        RECT 52.700 105.935 53.775 106.105 ;
        RECT 52.035 105.335 52.405 105.795 ;
        RECT 52.700 105.595 52.870 105.935 ;
        RECT 53.040 105.335 53.370 105.765 ;
        RECT 53.605 105.595 53.775 105.935 ;
        RECT 53.945 105.835 54.115 106.615 ;
        RECT 54.285 106.395 54.455 106.985 ;
        RECT 54.625 106.585 54.975 107.205 ;
        RECT 54.285 106.005 54.750 106.395 ;
        RECT 55.145 106.135 55.315 107.495 ;
        RECT 55.485 106.305 55.945 107.355 ;
        RECT 54.920 105.965 55.315 106.135 ;
        RECT 54.920 105.835 55.090 105.965 ;
        RECT 53.945 105.505 54.625 105.835 ;
        RECT 54.840 105.505 55.090 105.835 ;
        RECT 55.260 105.335 55.510 105.795 ;
        RECT 55.680 105.520 56.005 106.305 ;
        RECT 56.175 105.505 56.345 107.625 ;
        RECT 56.515 107.505 56.845 107.885 ;
        RECT 57.015 107.335 57.270 107.625 ;
        RECT 56.520 107.165 57.270 107.335 ;
        RECT 56.520 106.175 56.750 107.165 ;
        RECT 57.505 107.065 57.715 107.885 ;
        RECT 57.885 107.085 58.215 107.715 ;
        RECT 56.920 106.345 57.270 106.995 ;
        RECT 57.885 106.485 58.135 107.085 ;
        RECT 58.385 107.065 58.615 107.885 ;
        RECT 58.825 107.135 60.035 107.885 ;
        RECT 58.305 106.645 58.635 106.895 ;
        RECT 56.520 106.005 57.270 106.175 ;
        RECT 56.515 105.335 56.845 105.835 ;
        RECT 57.015 105.505 57.270 106.005 ;
        RECT 57.505 105.335 57.715 106.475 ;
        RECT 57.885 105.505 58.215 106.485 ;
        RECT 58.385 105.335 58.615 106.475 ;
        RECT 58.825 106.425 59.345 106.965 ;
        RECT 59.515 106.595 60.035 107.135 ;
        RECT 60.245 107.065 60.475 107.885 ;
        RECT 60.645 107.085 60.975 107.715 ;
        RECT 60.225 106.645 60.555 106.895 ;
        RECT 60.725 106.485 60.975 107.085 ;
        RECT 61.145 107.065 61.355 107.885 ;
        RECT 61.675 107.335 61.845 107.715 ;
        RECT 62.025 107.505 62.355 107.885 ;
        RECT 61.675 107.165 62.340 107.335 ;
        RECT 62.535 107.210 62.795 107.715 ;
        RECT 61.605 106.615 61.935 106.985 ;
        RECT 62.170 106.910 62.340 107.165 ;
        RECT 58.825 105.335 60.035 106.425 ;
        RECT 60.245 105.335 60.475 106.475 ;
        RECT 60.645 105.505 60.975 106.485 ;
        RECT 62.170 106.580 62.455 106.910 ;
        RECT 61.145 105.335 61.355 106.475 ;
        RECT 62.170 106.435 62.340 106.580 ;
        RECT 61.675 106.265 62.340 106.435 ;
        RECT 62.625 106.410 62.795 107.210 ;
        RECT 62.965 107.160 63.255 107.885 ;
        RECT 63.735 107.415 63.905 107.885 ;
        RECT 64.075 107.235 64.405 107.715 ;
        RECT 64.575 107.415 64.745 107.885 ;
        RECT 64.915 107.235 65.245 107.715 ;
        RECT 63.480 107.065 65.245 107.235 ;
        RECT 65.415 107.075 65.585 107.885 ;
        RECT 65.785 107.505 66.855 107.675 ;
        RECT 65.785 107.150 66.105 107.505 ;
        RECT 63.480 106.515 63.890 107.065 ;
        RECT 65.780 106.895 66.105 107.150 ;
        RECT 64.075 106.685 66.105 106.895 ;
        RECT 65.760 106.675 66.105 106.685 ;
        RECT 66.275 106.935 66.515 107.335 ;
        RECT 66.685 107.275 66.855 107.505 ;
        RECT 67.025 107.445 67.215 107.885 ;
        RECT 67.385 107.435 68.335 107.715 ;
        RECT 68.555 107.525 68.905 107.695 ;
        RECT 66.685 107.105 67.215 107.275 ;
        RECT 61.675 105.505 61.845 106.265 ;
        RECT 62.025 105.335 62.355 106.095 ;
        RECT 62.525 105.505 62.795 106.410 ;
        RECT 62.965 105.335 63.255 106.500 ;
        RECT 63.480 106.345 65.205 106.515 ;
        RECT 63.735 105.335 63.905 106.175 ;
        RECT 64.115 105.505 64.365 106.345 ;
        RECT 64.575 105.335 64.745 106.175 ;
        RECT 64.915 105.505 65.205 106.345 ;
        RECT 65.415 105.335 65.585 106.395 ;
        RECT 65.760 106.055 65.930 106.675 ;
        RECT 66.275 106.565 66.815 106.935 ;
        RECT 66.995 106.825 67.215 107.105 ;
        RECT 67.385 106.655 67.555 107.435 ;
        RECT 67.150 106.485 67.555 106.655 ;
        RECT 67.725 106.645 68.075 107.265 ;
        RECT 67.150 106.395 67.320 106.485 ;
        RECT 68.245 106.475 68.455 107.265 ;
        RECT 66.100 106.225 67.320 106.395 ;
        RECT 67.780 106.315 68.455 106.475 ;
        RECT 65.760 105.885 66.560 106.055 ;
        RECT 65.880 105.335 66.210 105.715 ;
        RECT 66.390 105.595 66.560 105.885 ;
        RECT 67.150 105.845 67.320 106.225 ;
        RECT 67.490 106.305 68.455 106.315 ;
        RECT 68.645 107.135 68.905 107.525 ;
        RECT 69.115 107.425 69.445 107.885 ;
        RECT 70.320 107.495 71.175 107.665 ;
        RECT 71.380 107.495 71.875 107.665 ;
        RECT 72.045 107.525 72.375 107.885 ;
        RECT 68.645 106.445 68.815 107.135 ;
        RECT 68.985 106.785 69.155 106.965 ;
        RECT 69.325 106.955 70.115 107.205 ;
        RECT 70.320 106.785 70.490 107.495 ;
        RECT 70.660 106.985 71.015 107.205 ;
        RECT 68.985 106.615 70.675 106.785 ;
        RECT 67.490 106.015 67.950 106.305 ;
        RECT 68.645 106.275 70.145 106.445 ;
        RECT 68.645 106.135 68.815 106.275 ;
        RECT 68.255 105.965 68.815 106.135 ;
        RECT 66.730 105.335 66.980 105.795 ;
        RECT 67.150 105.505 68.020 105.845 ;
        RECT 68.255 105.505 68.425 105.965 ;
        RECT 69.260 105.935 70.335 106.105 ;
        RECT 68.595 105.335 68.965 105.795 ;
        RECT 69.260 105.595 69.430 105.935 ;
        RECT 69.600 105.335 69.930 105.765 ;
        RECT 70.165 105.595 70.335 105.935 ;
        RECT 70.505 105.835 70.675 106.615 ;
        RECT 70.845 106.395 71.015 106.985 ;
        RECT 71.185 106.585 71.535 107.205 ;
        RECT 70.845 106.005 71.310 106.395 ;
        RECT 71.705 106.135 71.875 107.495 ;
        RECT 72.045 106.305 72.505 107.355 ;
        RECT 71.480 105.965 71.875 106.135 ;
        RECT 71.480 105.835 71.650 105.965 ;
        RECT 70.505 105.505 71.185 105.835 ;
        RECT 71.400 105.505 71.650 105.835 ;
        RECT 71.820 105.335 72.070 105.795 ;
        RECT 72.240 105.520 72.565 106.305 ;
        RECT 72.735 105.505 72.905 107.625 ;
        RECT 73.075 107.505 73.405 107.885 ;
        RECT 73.575 107.335 73.830 107.625 ;
        RECT 73.080 107.165 73.830 107.335 ;
        RECT 75.015 107.335 75.185 107.715 ;
        RECT 75.365 107.505 75.695 107.885 ;
        RECT 75.015 107.165 75.680 107.335 ;
        RECT 75.875 107.210 76.135 107.715 ;
        RECT 76.615 107.415 76.785 107.885 ;
        RECT 76.955 107.235 77.285 107.715 ;
        RECT 77.455 107.415 77.625 107.885 ;
        RECT 77.795 107.235 78.125 107.715 ;
        RECT 73.080 106.175 73.310 107.165 ;
        RECT 73.480 106.345 73.830 106.995 ;
        RECT 74.945 106.615 75.275 106.985 ;
        RECT 75.510 106.910 75.680 107.165 ;
        RECT 75.510 106.580 75.795 106.910 ;
        RECT 75.510 106.435 75.680 106.580 ;
        RECT 75.015 106.265 75.680 106.435 ;
        RECT 75.965 106.410 76.135 107.210 ;
        RECT 73.080 106.005 73.830 106.175 ;
        RECT 73.075 105.335 73.405 105.835 ;
        RECT 73.575 105.505 73.830 106.005 ;
        RECT 75.015 105.505 75.185 106.265 ;
        RECT 75.365 105.335 75.695 106.095 ;
        RECT 75.865 105.505 76.135 106.410 ;
        RECT 76.360 107.065 78.125 107.235 ;
        RECT 78.295 107.075 78.465 107.885 ;
        RECT 78.665 107.505 79.735 107.675 ;
        RECT 78.665 107.150 78.985 107.505 ;
        RECT 76.360 106.515 76.770 107.065 ;
        RECT 78.660 106.895 78.985 107.150 ;
        RECT 76.955 106.685 78.985 106.895 ;
        RECT 78.640 106.675 78.985 106.685 ;
        RECT 79.155 106.935 79.395 107.335 ;
        RECT 79.565 107.275 79.735 107.505 ;
        RECT 79.905 107.445 80.095 107.885 ;
        RECT 80.265 107.435 81.215 107.715 ;
        RECT 81.435 107.525 81.785 107.695 ;
        RECT 79.565 107.105 80.095 107.275 ;
        RECT 76.360 106.345 78.085 106.515 ;
        RECT 76.615 105.335 76.785 106.175 ;
        RECT 76.995 105.505 77.245 106.345 ;
        RECT 77.455 105.335 77.625 106.175 ;
        RECT 77.795 105.505 78.085 106.345 ;
        RECT 78.295 105.335 78.465 106.395 ;
        RECT 78.640 106.055 78.810 106.675 ;
        RECT 79.155 106.565 79.695 106.935 ;
        RECT 79.875 106.825 80.095 107.105 ;
        RECT 80.265 106.655 80.435 107.435 ;
        RECT 80.030 106.485 80.435 106.655 ;
        RECT 80.605 106.645 80.955 107.265 ;
        RECT 80.030 106.395 80.200 106.485 ;
        RECT 81.125 106.475 81.335 107.265 ;
        RECT 78.980 106.225 80.200 106.395 ;
        RECT 80.660 106.315 81.335 106.475 ;
        RECT 78.640 105.885 79.440 106.055 ;
        RECT 78.760 105.335 79.090 105.715 ;
        RECT 79.270 105.595 79.440 105.885 ;
        RECT 80.030 105.845 80.200 106.225 ;
        RECT 80.370 106.305 81.335 106.315 ;
        RECT 81.525 107.135 81.785 107.525 ;
        RECT 81.995 107.425 82.325 107.885 ;
        RECT 83.200 107.495 84.055 107.665 ;
        RECT 84.260 107.495 84.755 107.665 ;
        RECT 84.925 107.525 85.255 107.885 ;
        RECT 81.525 106.445 81.695 107.135 ;
        RECT 81.865 106.785 82.035 106.965 ;
        RECT 82.205 106.955 82.995 107.205 ;
        RECT 83.200 106.785 83.370 107.495 ;
        RECT 83.540 106.985 83.895 107.205 ;
        RECT 81.865 106.615 83.555 106.785 ;
        RECT 80.370 106.015 80.830 106.305 ;
        RECT 81.525 106.275 83.025 106.445 ;
        RECT 81.525 106.135 81.695 106.275 ;
        RECT 81.135 105.965 81.695 106.135 ;
        RECT 79.610 105.335 79.860 105.795 ;
        RECT 80.030 105.505 80.900 105.845 ;
        RECT 81.135 105.505 81.305 105.965 ;
        RECT 82.140 105.935 83.215 106.105 ;
        RECT 81.475 105.335 81.845 105.795 ;
        RECT 82.140 105.595 82.310 105.935 ;
        RECT 82.480 105.335 82.810 105.765 ;
        RECT 83.045 105.595 83.215 105.935 ;
        RECT 83.385 105.835 83.555 106.615 ;
        RECT 83.725 106.395 83.895 106.985 ;
        RECT 84.065 106.585 84.415 107.205 ;
        RECT 83.725 106.005 84.190 106.395 ;
        RECT 84.585 106.135 84.755 107.495 ;
        RECT 84.925 106.305 85.385 107.355 ;
        RECT 84.360 105.965 84.755 106.135 ;
        RECT 84.360 105.835 84.530 105.965 ;
        RECT 83.385 105.505 84.065 105.835 ;
        RECT 84.280 105.505 84.530 105.835 ;
        RECT 84.700 105.335 84.950 105.795 ;
        RECT 85.120 105.520 85.445 106.305 ;
        RECT 85.615 105.505 85.785 107.625 ;
        RECT 85.955 107.505 86.285 107.885 ;
        RECT 86.455 107.335 86.710 107.625 ;
        RECT 85.960 107.165 86.710 107.335 ;
        RECT 87.435 107.335 87.605 107.715 ;
        RECT 87.785 107.505 88.115 107.885 ;
        RECT 87.435 107.165 88.100 107.335 ;
        RECT 88.295 107.210 88.555 107.715 ;
        RECT 85.960 106.175 86.190 107.165 ;
        RECT 86.360 106.345 86.710 106.995 ;
        RECT 87.365 106.615 87.695 106.985 ;
        RECT 87.930 106.910 88.100 107.165 ;
        RECT 87.930 106.580 88.215 106.910 ;
        RECT 87.930 106.435 88.100 106.580 ;
        RECT 87.435 106.265 88.100 106.435 ;
        RECT 88.385 106.410 88.555 107.210 ;
        RECT 88.725 107.160 89.015 107.885 ;
        RECT 89.495 107.415 89.665 107.885 ;
        RECT 89.835 107.235 90.165 107.715 ;
        RECT 90.335 107.415 90.505 107.885 ;
        RECT 90.675 107.235 91.005 107.715 ;
        RECT 89.240 107.065 91.005 107.235 ;
        RECT 91.175 107.075 91.345 107.885 ;
        RECT 91.545 107.505 92.615 107.675 ;
        RECT 91.545 107.150 91.865 107.505 ;
        RECT 89.240 106.515 89.650 107.065 ;
        RECT 91.540 106.895 91.865 107.150 ;
        RECT 89.835 106.685 91.865 106.895 ;
        RECT 91.520 106.675 91.865 106.685 ;
        RECT 92.035 106.935 92.275 107.335 ;
        RECT 92.445 107.275 92.615 107.505 ;
        RECT 92.785 107.445 92.975 107.885 ;
        RECT 93.145 107.435 94.095 107.715 ;
        RECT 94.315 107.525 94.665 107.695 ;
        RECT 92.445 107.105 92.975 107.275 ;
        RECT 85.960 106.005 86.710 106.175 ;
        RECT 85.955 105.335 86.285 105.835 ;
        RECT 86.455 105.505 86.710 106.005 ;
        RECT 87.435 105.505 87.605 106.265 ;
        RECT 87.785 105.335 88.115 106.095 ;
        RECT 88.285 105.505 88.555 106.410 ;
        RECT 88.725 105.335 89.015 106.500 ;
        RECT 89.240 106.345 90.965 106.515 ;
        RECT 89.495 105.335 89.665 106.175 ;
        RECT 89.875 105.505 90.125 106.345 ;
        RECT 90.335 105.335 90.505 106.175 ;
        RECT 90.675 105.505 90.965 106.345 ;
        RECT 91.175 105.335 91.345 106.395 ;
        RECT 91.520 106.055 91.690 106.675 ;
        RECT 92.035 106.565 92.575 106.935 ;
        RECT 92.755 106.825 92.975 107.105 ;
        RECT 93.145 106.655 93.315 107.435 ;
        RECT 92.910 106.485 93.315 106.655 ;
        RECT 93.485 106.645 93.835 107.265 ;
        RECT 92.910 106.395 93.080 106.485 ;
        RECT 94.005 106.475 94.215 107.265 ;
        RECT 91.860 106.225 93.080 106.395 ;
        RECT 93.540 106.315 94.215 106.475 ;
        RECT 91.520 105.885 92.320 106.055 ;
        RECT 91.640 105.335 91.970 105.715 ;
        RECT 92.150 105.595 92.320 105.885 ;
        RECT 92.910 105.845 93.080 106.225 ;
        RECT 93.250 106.305 94.215 106.315 ;
        RECT 94.405 107.135 94.665 107.525 ;
        RECT 94.875 107.425 95.205 107.885 ;
        RECT 96.080 107.495 96.935 107.665 ;
        RECT 97.140 107.495 97.635 107.665 ;
        RECT 97.805 107.525 98.135 107.885 ;
        RECT 94.405 106.445 94.575 107.135 ;
        RECT 94.745 106.785 94.915 106.965 ;
        RECT 95.085 106.955 95.875 107.205 ;
        RECT 96.080 106.785 96.250 107.495 ;
        RECT 96.420 106.985 96.775 107.205 ;
        RECT 94.745 106.615 96.435 106.785 ;
        RECT 93.250 106.015 93.710 106.305 ;
        RECT 94.405 106.275 95.905 106.445 ;
        RECT 94.405 106.135 94.575 106.275 ;
        RECT 94.015 105.965 94.575 106.135 ;
        RECT 92.490 105.335 92.740 105.795 ;
        RECT 92.910 105.505 93.780 105.845 ;
        RECT 94.015 105.505 94.185 105.965 ;
        RECT 95.020 105.935 96.095 106.105 ;
        RECT 94.355 105.335 94.725 105.795 ;
        RECT 95.020 105.595 95.190 105.935 ;
        RECT 95.360 105.335 95.690 105.765 ;
        RECT 95.925 105.595 96.095 105.935 ;
        RECT 96.265 105.835 96.435 106.615 ;
        RECT 96.605 106.395 96.775 106.985 ;
        RECT 96.945 106.585 97.295 107.205 ;
        RECT 96.605 106.005 97.070 106.395 ;
        RECT 97.465 106.135 97.635 107.495 ;
        RECT 97.805 106.305 98.265 107.355 ;
        RECT 97.240 105.965 97.635 106.135 ;
        RECT 97.240 105.835 97.410 105.965 ;
        RECT 96.265 105.505 96.945 105.835 ;
        RECT 97.160 105.505 97.410 105.835 ;
        RECT 97.580 105.335 97.830 105.795 ;
        RECT 98.000 105.520 98.325 106.305 ;
        RECT 98.495 105.505 98.665 107.625 ;
        RECT 98.835 107.505 99.165 107.885 ;
        RECT 99.335 107.335 99.590 107.625 ;
        RECT 98.840 107.165 99.590 107.335 ;
        RECT 98.840 106.175 99.070 107.165 ;
        RECT 99.825 107.065 100.035 107.885 ;
        RECT 100.205 107.085 100.535 107.715 ;
        RECT 99.240 106.345 99.590 106.995 ;
        RECT 100.205 106.485 100.455 107.085 ;
        RECT 100.705 107.065 100.935 107.885 ;
        RECT 101.145 107.135 102.355 107.885 ;
        RECT 100.625 106.645 100.955 106.895 ;
        RECT 98.840 106.005 99.590 106.175 ;
        RECT 98.835 105.335 99.165 105.835 ;
        RECT 99.335 105.505 99.590 106.005 ;
        RECT 99.825 105.335 100.035 106.475 ;
        RECT 100.205 105.505 100.535 106.485 ;
        RECT 100.705 105.335 100.935 106.475 ;
        RECT 101.145 106.425 101.665 106.965 ;
        RECT 101.835 106.595 102.355 107.135 ;
        RECT 102.565 107.065 102.795 107.885 ;
        RECT 102.965 107.085 103.295 107.715 ;
        RECT 102.545 106.645 102.875 106.895 ;
        RECT 103.045 106.485 103.295 107.085 ;
        RECT 103.465 107.065 103.675 107.885 ;
        RECT 104.215 107.415 104.385 107.885 ;
        RECT 104.555 107.235 104.885 107.715 ;
        RECT 105.055 107.415 105.225 107.885 ;
        RECT 105.395 107.235 105.725 107.715 ;
        RECT 103.960 107.065 105.725 107.235 ;
        RECT 105.895 107.075 106.065 107.885 ;
        RECT 106.265 107.505 107.335 107.675 ;
        RECT 106.265 107.150 106.585 107.505 ;
        RECT 101.145 105.335 102.355 106.425 ;
        RECT 102.565 105.335 102.795 106.475 ;
        RECT 102.965 105.505 103.295 106.485 ;
        RECT 103.960 106.515 104.370 107.065 ;
        RECT 106.260 106.895 106.585 107.150 ;
        RECT 104.555 106.685 106.585 106.895 ;
        RECT 106.240 106.675 106.585 106.685 ;
        RECT 106.755 106.935 106.995 107.335 ;
        RECT 107.165 107.275 107.335 107.505 ;
        RECT 107.505 107.445 107.695 107.885 ;
        RECT 107.865 107.435 108.815 107.715 ;
        RECT 109.035 107.525 109.385 107.695 ;
        RECT 107.165 107.105 107.695 107.275 ;
        RECT 103.465 105.335 103.675 106.475 ;
        RECT 103.960 106.345 105.685 106.515 ;
        RECT 104.215 105.335 104.385 106.175 ;
        RECT 104.595 105.505 104.845 106.345 ;
        RECT 105.055 105.335 105.225 106.175 ;
        RECT 105.395 105.505 105.685 106.345 ;
        RECT 105.895 105.335 106.065 106.395 ;
        RECT 106.240 106.055 106.410 106.675 ;
        RECT 106.755 106.565 107.295 106.935 ;
        RECT 107.475 106.825 107.695 107.105 ;
        RECT 107.865 106.655 108.035 107.435 ;
        RECT 107.630 106.485 108.035 106.655 ;
        RECT 108.205 106.645 108.555 107.265 ;
        RECT 107.630 106.395 107.800 106.485 ;
        RECT 108.725 106.475 108.935 107.265 ;
        RECT 106.580 106.225 107.800 106.395 ;
        RECT 108.260 106.315 108.935 106.475 ;
        RECT 106.240 105.885 107.040 106.055 ;
        RECT 106.360 105.335 106.690 105.715 ;
        RECT 106.870 105.595 107.040 105.885 ;
        RECT 107.630 105.845 107.800 106.225 ;
        RECT 107.970 106.305 108.935 106.315 ;
        RECT 109.125 107.135 109.385 107.525 ;
        RECT 109.595 107.425 109.925 107.885 ;
        RECT 110.800 107.495 111.655 107.665 ;
        RECT 111.860 107.495 112.355 107.665 ;
        RECT 112.525 107.525 112.855 107.885 ;
        RECT 109.125 106.445 109.295 107.135 ;
        RECT 109.465 106.785 109.635 106.965 ;
        RECT 109.805 106.955 110.595 107.205 ;
        RECT 110.800 106.785 110.970 107.495 ;
        RECT 111.140 106.985 111.495 107.205 ;
        RECT 109.465 106.615 111.155 106.785 ;
        RECT 107.970 106.015 108.430 106.305 ;
        RECT 109.125 106.275 110.625 106.445 ;
        RECT 109.125 106.135 109.295 106.275 ;
        RECT 108.735 105.965 109.295 106.135 ;
        RECT 107.210 105.335 107.460 105.795 ;
        RECT 107.630 105.505 108.500 105.845 ;
        RECT 108.735 105.505 108.905 105.965 ;
        RECT 109.740 105.935 110.815 106.105 ;
        RECT 109.075 105.335 109.445 105.795 ;
        RECT 109.740 105.595 109.910 105.935 ;
        RECT 110.080 105.335 110.410 105.765 ;
        RECT 110.645 105.595 110.815 105.935 ;
        RECT 110.985 105.835 111.155 106.615 ;
        RECT 111.325 106.395 111.495 106.985 ;
        RECT 111.665 106.585 112.015 107.205 ;
        RECT 111.325 106.005 111.790 106.395 ;
        RECT 112.185 106.135 112.355 107.495 ;
        RECT 112.525 106.305 112.985 107.355 ;
        RECT 111.960 105.965 112.355 106.135 ;
        RECT 111.960 105.835 112.130 105.965 ;
        RECT 110.985 105.505 111.665 105.835 ;
        RECT 111.880 105.505 112.130 105.835 ;
        RECT 112.300 105.335 112.550 105.795 ;
        RECT 112.720 105.520 113.045 106.305 ;
        RECT 113.215 105.505 113.385 107.625 ;
        RECT 113.555 107.505 113.885 107.885 ;
        RECT 114.055 107.335 114.310 107.625 ;
        RECT 113.560 107.165 114.310 107.335 ;
        RECT 113.560 106.175 113.790 107.165 ;
        RECT 114.485 107.160 114.775 107.885 ;
        RECT 115.870 107.335 116.125 107.625 ;
        RECT 116.295 107.505 116.625 107.885 ;
        RECT 115.870 107.165 116.620 107.335 ;
        RECT 113.960 106.345 114.310 106.995 ;
        RECT 113.560 106.005 114.310 106.175 ;
        RECT 113.555 105.335 113.885 105.835 ;
        RECT 114.055 105.505 114.310 106.005 ;
        RECT 114.485 105.335 114.775 106.500 ;
        RECT 115.870 106.345 116.220 106.995 ;
        RECT 116.390 106.175 116.620 107.165 ;
        RECT 115.870 106.005 116.620 106.175 ;
        RECT 115.870 105.505 116.125 106.005 ;
        RECT 116.295 105.335 116.625 105.835 ;
        RECT 116.795 105.505 116.965 107.625 ;
        RECT 117.325 107.525 117.655 107.885 ;
        RECT 117.825 107.495 118.320 107.665 ;
        RECT 118.525 107.495 119.380 107.665 ;
        RECT 117.195 106.305 117.655 107.355 ;
        RECT 117.135 105.520 117.460 106.305 ;
        RECT 117.825 106.135 117.995 107.495 ;
        RECT 118.165 106.585 118.515 107.205 ;
        RECT 118.685 106.985 119.040 107.205 ;
        RECT 118.685 106.395 118.855 106.985 ;
        RECT 119.210 106.785 119.380 107.495 ;
        RECT 120.255 107.425 120.585 107.885 ;
        RECT 120.795 107.525 121.145 107.695 ;
        RECT 119.585 106.955 120.375 107.205 ;
        RECT 120.795 107.135 121.055 107.525 ;
        RECT 121.365 107.435 122.315 107.715 ;
        RECT 122.485 107.445 122.675 107.885 ;
        RECT 122.845 107.505 123.915 107.675 ;
        RECT 120.545 106.785 120.715 106.965 ;
        RECT 117.825 105.965 118.220 106.135 ;
        RECT 118.390 106.005 118.855 106.395 ;
        RECT 119.025 106.615 120.715 106.785 ;
        RECT 118.050 105.835 118.220 105.965 ;
        RECT 119.025 105.835 119.195 106.615 ;
        RECT 120.885 106.445 121.055 107.135 ;
        RECT 119.555 106.275 121.055 106.445 ;
        RECT 121.245 106.475 121.455 107.265 ;
        RECT 121.625 106.645 121.975 107.265 ;
        RECT 122.145 106.655 122.315 107.435 ;
        RECT 122.845 107.275 123.015 107.505 ;
        RECT 122.485 107.105 123.015 107.275 ;
        RECT 122.485 106.825 122.705 107.105 ;
        RECT 123.185 106.935 123.425 107.335 ;
        RECT 122.145 106.485 122.550 106.655 ;
        RECT 122.885 106.565 123.425 106.935 ;
        RECT 123.595 107.150 123.915 107.505 ;
        RECT 123.595 106.895 123.920 107.150 ;
        RECT 124.115 107.075 124.285 107.885 ;
        RECT 124.455 107.235 124.785 107.715 ;
        RECT 124.955 107.415 125.125 107.885 ;
        RECT 125.295 107.235 125.625 107.715 ;
        RECT 125.795 107.415 125.965 107.885 ;
        RECT 124.455 107.065 126.220 107.235 ;
        RECT 126.445 107.135 127.655 107.885 ;
        RECT 123.595 106.685 125.625 106.895 ;
        RECT 123.595 106.675 123.940 106.685 ;
        RECT 121.245 106.315 121.920 106.475 ;
        RECT 122.380 106.395 122.550 106.485 ;
        RECT 121.245 106.305 122.210 106.315 ;
        RECT 120.885 106.135 121.055 106.275 ;
        RECT 117.630 105.335 117.880 105.795 ;
        RECT 118.050 105.505 118.300 105.835 ;
        RECT 118.515 105.505 119.195 105.835 ;
        RECT 119.365 105.935 120.440 106.105 ;
        RECT 120.885 105.965 121.445 106.135 ;
        RECT 121.750 106.015 122.210 106.305 ;
        RECT 122.380 106.225 123.600 106.395 ;
        RECT 119.365 105.595 119.535 105.935 ;
        RECT 119.770 105.335 120.100 105.765 ;
        RECT 120.270 105.595 120.440 105.935 ;
        RECT 120.735 105.335 121.105 105.795 ;
        RECT 121.275 105.505 121.445 105.965 ;
        RECT 122.380 105.845 122.550 106.225 ;
        RECT 123.770 106.055 123.940 106.675 ;
        RECT 125.810 106.515 126.220 107.065 ;
        RECT 121.680 105.505 122.550 105.845 ;
        RECT 123.140 105.885 123.940 106.055 ;
        RECT 122.720 105.335 122.970 105.795 ;
        RECT 123.140 105.595 123.310 105.885 ;
        RECT 123.490 105.335 123.820 105.715 ;
        RECT 124.115 105.335 124.285 106.395 ;
        RECT 124.495 106.345 126.220 106.515 ;
        RECT 126.445 106.425 126.965 106.965 ;
        RECT 127.135 106.595 127.655 107.135 ;
        RECT 124.495 105.505 124.785 106.345 ;
        RECT 124.955 105.335 125.125 106.175 ;
        RECT 125.335 105.505 125.585 106.345 ;
        RECT 125.795 105.335 125.965 106.175 ;
        RECT 126.445 105.335 127.655 106.425 ;
        RECT 14.580 105.165 127.740 105.335 ;
        RECT 14.665 104.075 15.875 105.165 ;
        RECT 14.665 103.365 15.185 103.905 ;
        RECT 15.355 103.535 15.875 104.075 ;
        RECT 16.045 104.075 18.635 105.165 ;
        RECT 18.810 104.730 24.155 105.165 ;
        RECT 16.045 103.555 17.255 104.075 ;
        RECT 17.425 103.385 18.635 103.905 ;
        RECT 20.400 103.480 20.750 104.730 ;
        RECT 24.325 104.000 24.615 105.165 ;
        RECT 24.785 104.075 27.375 105.165 ;
        RECT 14.665 102.615 15.875 103.365 ;
        RECT 16.045 102.615 18.635 103.385 ;
        RECT 22.230 103.160 22.570 103.990 ;
        RECT 24.785 103.555 25.995 104.075 ;
        RECT 27.585 104.025 27.815 105.165 ;
        RECT 27.985 104.015 28.315 104.995 ;
        RECT 28.485 104.025 28.695 105.165 ;
        RECT 28.930 104.495 29.185 104.995 ;
        RECT 29.355 104.665 29.685 105.165 ;
        RECT 28.930 104.325 29.680 104.495 ;
        RECT 26.165 103.385 27.375 103.905 ;
        RECT 27.565 103.605 27.895 103.855 ;
        RECT 18.810 102.615 24.155 103.160 ;
        RECT 24.325 102.615 24.615 103.340 ;
        RECT 24.785 102.615 27.375 103.385 ;
        RECT 27.585 102.615 27.815 103.435 ;
        RECT 28.065 103.415 28.315 104.015 ;
        RECT 28.930 103.505 29.280 104.155 ;
        RECT 27.985 102.785 28.315 103.415 ;
        RECT 28.485 102.615 28.695 103.435 ;
        RECT 29.450 103.335 29.680 104.325 ;
        RECT 28.930 103.165 29.680 103.335 ;
        RECT 28.930 102.875 29.185 103.165 ;
        RECT 29.355 102.615 29.685 102.995 ;
        RECT 29.855 102.875 30.025 104.995 ;
        RECT 30.195 104.195 30.520 104.980 ;
        RECT 30.690 104.705 30.940 105.165 ;
        RECT 31.110 104.665 31.360 104.995 ;
        RECT 31.575 104.665 32.255 104.995 ;
        RECT 31.110 104.535 31.280 104.665 ;
        RECT 30.885 104.365 31.280 104.535 ;
        RECT 30.255 103.145 30.715 104.195 ;
        RECT 30.885 103.005 31.055 104.365 ;
        RECT 31.450 104.105 31.915 104.495 ;
        RECT 31.225 103.295 31.575 103.915 ;
        RECT 31.745 103.515 31.915 104.105 ;
        RECT 32.085 103.885 32.255 104.665 ;
        RECT 32.425 104.565 32.595 104.905 ;
        RECT 32.830 104.735 33.160 105.165 ;
        RECT 33.330 104.565 33.500 104.905 ;
        RECT 33.795 104.705 34.165 105.165 ;
        RECT 32.425 104.395 33.500 104.565 ;
        RECT 34.335 104.535 34.505 104.995 ;
        RECT 34.740 104.655 35.610 104.995 ;
        RECT 35.780 104.705 36.030 105.165 ;
        RECT 33.945 104.365 34.505 104.535 ;
        RECT 33.945 104.225 34.115 104.365 ;
        RECT 32.615 104.055 34.115 104.225 ;
        RECT 34.810 104.195 35.270 104.485 ;
        RECT 32.085 103.715 33.775 103.885 ;
        RECT 31.745 103.295 32.100 103.515 ;
        RECT 32.270 103.005 32.440 103.715 ;
        RECT 32.645 103.295 33.435 103.545 ;
        RECT 33.605 103.535 33.775 103.715 ;
        RECT 33.945 103.365 34.115 104.055 ;
        RECT 30.385 102.615 30.715 102.975 ;
        RECT 30.885 102.835 31.380 103.005 ;
        RECT 31.585 102.835 32.440 103.005 ;
        RECT 33.315 102.615 33.645 103.075 ;
        RECT 33.855 102.975 34.115 103.365 ;
        RECT 34.305 104.185 35.270 104.195 ;
        RECT 35.440 104.275 35.610 104.655 ;
        RECT 36.200 104.615 36.370 104.905 ;
        RECT 36.550 104.785 36.880 105.165 ;
        RECT 36.200 104.445 37.000 104.615 ;
        RECT 34.305 104.025 34.980 104.185 ;
        RECT 35.440 104.105 36.660 104.275 ;
        RECT 34.305 103.235 34.515 104.025 ;
        RECT 35.440 104.015 35.610 104.105 ;
        RECT 34.685 103.235 35.035 103.855 ;
        RECT 35.205 103.845 35.610 104.015 ;
        RECT 35.205 103.065 35.375 103.845 ;
        RECT 35.545 103.395 35.765 103.675 ;
        RECT 35.945 103.565 36.485 103.935 ;
        RECT 36.830 103.825 37.000 104.445 ;
        RECT 37.175 104.105 37.345 105.165 ;
        RECT 37.555 104.155 37.845 104.995 ;
        RECT 38.015 104.325 38.185 105.165 ;
        RECT 38.395 104.155 38.645 104.995 ;
        RECT 38.855 104.325 39.025 105.165 ;
        RECT 39.815 104.325 39.985 105.165 ;
        RECT 40.195 104.155 40.445 104.995 ;
        RECT 40.655 104.325 40.825 105.165 ;
        RECT 40.995 104.155 41.285 104.995 ;
        RECT 37.555 103.985 39.280 104.155 ;
        RECT 35.545 103.225 36.075 103.395 ;
        RECT 33.855 102.805 34.205 102.975 ;
        RECT 34.425 102.785 35.375 103.065 ;
        RECT 35.545 102.615 35.735 103.055 ;
        RECT 35.905 102.995 36.075 103.225 ;
        RECT 36.245 103.165 36.485 103.565 ;
        RECT 36.655 103.815 37.000 103.825 ;
        RECT 36.655 103.605 38.685 103.815 ;
        RECT 36.655 103.350 36.980 103.605 ;
        RECT 38.870 103.435 39.280 103.985 ;
        RECT 36.655 102.995 36.975 103.350 ;
        RECT 35.905 102.825 36.975 102.995 ;
        RECT 37.175 102.615 37.345 103.425 ;
        RECT 37.515 103.265 39.280 103.435 ;
        RECT 39.560 103.985 41.285 104.155 ;
        RECT 41.495 104.105 41.665 105.165 ;
        RECT 41.960 104.785 42.290 105.165 ;
        RECT 42.470 104.615 42.640 104.905 ;
        RECT 42.810 104.705 43.060 105.165 ;
        RECT 41.840 104.445 42.640 104.615 ;
        RECT 43.230 104.655 44.100 104.995 ;
        RECT 39.560 103.435 39.970 103.985 ;
        RECT 41.840 103.825 42.010 104.445 ;
        RECT 43.230 104.275 43.400 104.655 ;
        RECT 44.335 104.535 44.505 104.995 ;
        RECT 44.675 104.705 45.045 105.165 ;
        RECT 45.340 104.565 45.510 104.905 ;
        RECT 45.680 104.735 46.010 105.165 ;
        RECT 46.245 104.565 46.415 104.905 ;
        RECT 42.180 104.105 43.400 104.275 ;
        RECT 43.570 104.195 44.030 104.485 ;
        RECT 44.335 104.365 44.895 104.535 ;
        RECT 45.340 104.395 46.415 104.565 ;
        RECT 46.585 104.665 47.265 104.995 ;
        RECT 47.480 104.665 47.730 104.995 ;
        RECT 47.900 104.705 48.150 105.165 ;
        RECT 44.725 104.225 44.895 104.365 ;
        RECT 43.570 104.185 44.535 104.195 ;
        RECT 43.230 104.015 43.400 104.105 ;
        RECT 43.860 104.025 44.535 104.185 ;
        RECT 41.840 103.815 42.185 103.825 ;
        RECT 40.155 103.605 42.185 103.815 ;
        RECT 39.560 103.265 41.325 103.435 ;
        RECT 37.515 102.785 37.845 103.265 ;
        RECT 38.015 102.615 38.185 103.085 ;
        RECT 38.355 102.785 38.685 103.265 ;
        RECT 38.855 102.615 39.025 103.085 ;
        RECT 39.815 102.615 39.985 103.085 ;
        RECT 40.155 102.785 40.485 103.265 ;
        RECT 40.655 102.615 40.825 103.085 ;
        RECT 40.995 102.785 41.325 103.265 ;
        RECT 41.495 102.615 41.665 103.425 ;
        RECT 41.860 103.350 42.185 103.605 ;
        RECT 41.865 102.995 42.185 103.350 ;
        RECT 42.355 103.565 42.895 103.935 ;
        RECT 43.230 103.845 43.635 104.015 ;
        RECT 42.355 103.165 42.595 103.565 ;
        RECT 43.075 103.395 43.295 103.675 ;
        RECT 42.765 103.225 43.295 103.395 ;
        RECT 42.765 102.995 42.935 103.225 ;
        RECT 43.465 103.065 43.635 103.845 ;
        RECT 43.805 103.235 44.155 103.855 ;
        RECT 44.325 103.235 44.535 104.025 ;
        RECT 44.725 104.055 46.225 104.225 ;
        RECT 44.725 103.365 44.895 104.055 ;
        RECT 46.585 103.885 46.755 104.665 ;
        RECT 47.560 104.535 47.730 104.665 ;
        RECT 45.065 103.715 46.755 103.885 ;
        RECT 46.925 104.105 47.390 104.495 ;
        RECT 47.560 104.365 47.955 104.535 ;
        RECT 45.065 103.535 45.235 103.715 ;
        RECT 41.865 102.825 42.935 102.995 ;
        RECT 43.105 102.615 43.295 103.055 ;
        RECT 43.465 102.785 44.415 103.065 ;
        RECT 44.725 102.975 44.985 103.365 ;
        RECT 45.405 103.295 46.195 103.545 ;
        RECT 44.635 102.805 44.985 102.975 ;
        RECT 45.195 102.615 45.525 103.075 ;
        RECT 46.400 103.005 46.570 103.715 ;
        RECT 46.925 103.515 47.095 104.105 ;
        RECT 46.740 103.295 47.095 103.515 ;
        RECT 47.265 103.295 47.615 103.915 ;
        RECT 47.785 103.005 47.955 104.365 ;
        RECT 48.320 104.195 48.645 104.980 ;
        RECT 48.125 103.145 48.585 104.195 ;
        RECT 46.400 102.835 47.255 103.005 ;
        RECT 47.460 102.835 47.955 103.005 ;
        RECT 48.125 102.615 48.455 102.975 ;
        RECT 48.815 102.875 48.985 104.995 ;
        RECT 49.155 104.665 49.485 105.165 ;
        RECT 49.655 104.495 49.910 104.995 ;
        RECT 49.160 104.325 49.910 104.495 ;
        RECT 49.160 103.335 49.390 104.325 ;
        RECT 49.560 103.505 49.910 104.155 ;
        RECT 50.085 104.000 50.375 105.165 ;
        RECT 51.525 104.025 51.735 105.165 ;
        RECT 51.905 104.015 52.235 104.995 ;
        RECT 52.405 104.025 52.635 105.165 ;
        RECT 53.155 104.325 53.325 105.165 ;
        RECT 53.535 104.155 53.785 104.995 ;
        RECT 53.995 104.325 54.165 105.165 ;
        RECT 54.335 104.155 54.625 104.995 ;
        RECT 49.160 103.165 49.910 103.335 ;
        RECT 49.155 102.615 49.485 102.995 ;
        RECT 49.655 102.875 49.910 103.165 ;
        RECT 50.085 102.615 50.375 103.340 ;
        RECT 51.525 102.615 51.735 103.435 ;
        RECT 51.905 103.415 52.155 104.015 ;
        RECT 52.900 103.985 54.625 104.155 ;
        RECT 54.835 104.105 55.005 105.165 ;
        RECT 55.300 104.785 55.630 105.165 ;
        RECT 55.810 104.615 55.980 104.905 ;
        RECT 56.150 104.705 56.400 105.165 ;
        RECT 55.180 104.445 55.980 104.615 ;
        RECT 56.570 104.655 57.440 104.995 ;
        RECT 52.325 103.605 52.655 103.855 ;
        RECT 52.900 103.435 53.310 103.985 ;
        RECT 55.180 103.825 55.350 104.445 ;
        RECT 56.570 104.275 56.740 104.655 ;
        RECT 57.675 104.535 57.845 104.995 ;
        RECT 58.015 104.705 58.385 105.165 ;
        RECT 58.680 104.565 58.850 104.905 ;
        RECT 59.020 104.735 59.350 105.165 ;
        RECT 59.585 104.565 59.755 104.905 ;
        RECT 55.520 104.105 56.740 104.275 ;
        RECT 56.910 104.195 57.370 104.485 ;
        RECT 57.675 104.365 58.235 104.535 ;
        RECT 58.680 104.395 59.755 104.565 ;
        RECT 59.925 104.665 60.605 104.995 ;
        RECT 60.820 104.665 61.070 104.995 ;
        RECT 61.240 104.705 61.490 105.165 ;
        RECT 58.065 104.225 58.235 104.365 ;
        RECT 56.910 104.185 57.875 104.195 ;
        RECT 56.570 104.015 56.740 104.105 ;
        RECT 57.200 104.025 57.875 104.185 ;
        RECT 55.180 103.815 55.525 103.825 ;
        RECT 53.495 103.605 55.525 103.815 ;
        RECT 51.905 102.785 52.235 103.415 ;
        RECT 52.405 102.615 52.635 103.435 ;
        RECT 52.900 103.265 54.665 103.435 ;
        RECT 53.155 102.615 53.325 103.085 ;
        RECT 53.495 102.785 53.825 103.265 ;
        RECT 53.995 102.615 54.165 103.085 ;
        RECT 54.335 102.785 54.665 103.265 ;
        RECT 54.835 102.615 55.005 103.425 ;
        RECT 55.200 103.350 55.525 103.605 ;
        RECT 55.205 102.995 55.525 103.350 ;
        RECT 55.695 103.565 56.235 103.935 ;
        RECT 56.570 103.845 56.975 104.015 ;
        RECT 55.695 103.165 55.935 103.565 ;
        RECT 56.415 103.395 56.635 103.675 ;
        RECT 56.105 103.225 56.635 103.395 ;
        RECT 56.105 102.995 56.275 103.225 ;
        RECT 56.805 103.065 56.975 103.845 ;
        RECT 57.145 103.235 57.495 103.855 ;
        RECT 57.665 103.235 57.875 104.025 ;
        RECT 58.065 104.055 59.565 104.225 ;
        RECT 58.065 103.365 58.235 104.055 ;
        RECT 59.925 103.885 60.095 104.665 ;
        RECT 60.900 104.535 61.070 104.665 ;
        RECT 58.405 103.715 60.095 103.885 ;
        RECT 60.265 104.105 60.730 104.495 ;
        RECT 60.900 104.365 61.295 104.535 ;
        RECT 58.405 103.535 58.575 103.715 ;
        RECT 55.205 102.825 56.275 102.995 ;
        RECT 56.445 102.615 56.635 103.055 ;
        RECT 56.805 102.785 57.755 103.065 ;
        RECT 58.065 102.975 58.325 103.365 ;
        RECT 58.745 103.295 59.535 103.545 ;
        RECT 57.975 102.805 58.325 102.975 ;
        RECT 58.535 102.615 58.865 103.075 ;
        RECT 59.740 103.005 59.910 103.715 ;
        RECT 60.265 103.515 60.435 104.105 ;
        RECT 60.080 103.295 60.435 103.515 ;
        RECT 60.605 103.295 60.955 103.915 ;
        RECT 61.125 103.005 61.295 104.365 ;
        RECT 61.660 104.195 61.985 104.980 ;
        RECT 61.465 103.145 61.925 104.195 ;
        RECT 59.740 102.835 60.595 103.005 ;
        RECT 60.800 102.835 61.295 103.005 ;
        RECT 61.465 102.615 61.795 102.975 ;
        RECT 62.155 102.875 62.325 104.995 ;
        RECT 62.495 104.665 62.825 105.165 ;
        RECT 62.995 104.495 63.250 104.995 ;
        RECT 62.500 104.325 63.250 104.495 ;
        RECT 63.735 104.325 63.905 105.165 ;
        RECT 62.500 103.335 62.730 104.325 ;
        RECT 64.115 104.155 64.365 104.995 ;
        RECT 64.575 104.325 64.745 105.165 ;
        RECT 64.915 104.155 65.205 104.995 ;
        RECT 62.900 103.505 63.250 104.155 ;
        RECT 63.480 103.985 65.205 104.155 ;
        RECT 65.415 104.105 65.585 105.165 ;
        RECT 65.880 104.785 66.210 105.165 ;
        RECT 66.390 104.615 66.560 104.905 ;
        RECT 66.730 104.705 66.980 105.165 ;
        RECT 65.760 104.445 66.560 104.615 ;
        RECT 67.150 104.655 68.020 104.995 ;
        RECT 63.480 103.435 63.890 103.985 ;
        RECT 65.760 103.825 65.930 104.445 ;
        RECT 67.150 104.275 67.320 104.655 ;
        RECT 68.255 104.535 68.425 104.995 ;
        RECT 68.595 104.705 68.965 105.165 ;
        RECT 69.260 104.565 69.430 104.905 ;
        RECT 69.600 104.735 69.930 105.165 ;
        RECT 70.165 104.565 70.335 104.905 ;
        RECT 66.100 104.105 67.320 104.275 ;
        RECT 67.490 104.195 67.950 104.485 ;
        RECT 68.255 104.365 68.815 104.535 ;
        RECT 69.260 104.395 70.335 104.565 ;
        RECT 70.505 104.665 71.185 104.995 ;
        RECT 71.400 104.665 71.650 104.995 ;
        RECT 71.820 104.705 72.070 105.165 ;
        RECT 68.645 104.225 68.815 104.365 ;
        RECT 67.490 104.185 68.455 104.195 ;
        RECT 67.150 104.015 67.320 104.105 ;
        RECT 67.780 104.025 68.455 104.185 ;
        RECT 65.760 103.815 66.105 103.825 ;
        RECT 64.075 103.605 66.105 103.815 ;
        RECT 62.500 103.165 63.250 103.335 ;
        RECT 63.480 103.265 65.245 103.435 ;
        RECT 62.495 102.615 62.825 102.995 ;
        RECT 62.995 102.875 63.250 103.165 ;
        RECT 63.735 102.615 63.905 103.085 ;
        RECT 64.075 102.785 64.405 103.265 ;
        RECT 64.575 102.615 64.745 103.085 ;
        RECT 64.915 102.785 65.245 103.265 ;
        RECT 65.415 102.615 65.585 103.425 ;
        RECT 65.780 103.350 66.105 103.605 ;
        RECT 65.785 102.995 66.105 103.350 ;
        RECT 66.275 103.565 66.815 103.935 ;
        RECT 67.150 103.845 67.555 104.015 ;
        RECT 66.275 103.165 66.515 103.565 ;
        RECT 66.995 103.395 67.215 103.675 ;
        RECT 66.685 103.225 67.215 103.395 ;
        RECT 66.685 102.995 66.855 103.225 ;
        RECT 67.385 103.065 67.555 103.845 ;
        RECT 67.725 103.235 68.075 103.855 ;
        RECT 68.245 103.235 68.455 104.025 ;
        RECT 68.645 104.055 70.145 104.225 ;
        RECT 68.645 103.365 68.815 104.055 ;
        RECT 70.505 103.885 70.675 104.665 ;
        RECT 71.480 104.535 71.650 104.665 ;
        RECT 68.985 103.715 70.675 103.885 ;
        RECT 70.845 104.105 71.310 104.495 ;
        RECT 71.480 104.365 71.875 104.535 ;
        RECT 68.985 103.535 69.155 103.715 ;
        RECT 65.785 102.825 66.855 102.995 ;
        RECT 67.025 102.615 67.215 103.055 ;
        RECT 67.385 102.785 68.335 103.065 ;
        RECT 68.645 102.975 68.905 103.365 ;
        RECT 69.325 103.295 70.115 103.545 ;
        RECT 68.555 102.805 68.905 102.975 ;
        RECT 69.115 102.615 69.445 103.075 ;
        RECT 70.320 103.005 70.490 103.715 ;
        RECT 70.845 103.515 71.015 104.105 ;
        RECT 70.660 103.295 71.015 103.515 ;
        RECT 71.185 103.295 71.535 103.915 ;
        RECT 71.705 103.005 71.875 104.365 ;
        RECT 72.240 104.195 72.565 104.980 ;
        RECT 72.045 103.145 72.505 104.195 ;
        RECT 70.320 102.835 71.175 103.005 ;
        RECT 71.380 102.835 71.875 103.005 ;
        RECT 72.045 102.615 72.375 102.975 ;
        RECT 72.735 102.875 72.905 104.995 ;
        RECT 73.075 104.665 73.405 105.165 ;
        RECT 73.575 104.495 73.830 104.995 ;
        RECT 73.080 104.325 73.830 104.495 ;
        RECT 73.080 103.335 73.310 104.325 ;
        RECT 73.480 103.505 73.830 104.155 ;
        RECT 74.005 104.075 75.675 105.165 ;
        RECT 74.005 103.555 74.755 104.075 ;
        RECT 75.845 104.000 76.135 105.165 ;
        RECT 76.615 104.325 76.785 105.165 ;
        RECT 76.995 104.155 77.245 104.995 ;
        RECT 77.455 104.325 77.625 105.165 ;
        RECT 77.795 104.155 78.085 104.995 ;
        RECT 76.360 103.985 78.085 104.155 ;
        RECT 78.295 104.105 78.465 105.165 ;
        RECT 78.760 104.785 79.090 105.165 ;
        RECT 79.270 104.615 79.440 104.905 ;
        RECT 79.610 104.705 79.860 105.165 ;
        RECT 78.640 104.445 79.440 104.615 ;
        RECT 80.030 104.655 80.900 104.995 ;
        RECT 74.925 103.385 75.675 103.905 ;
        RECT 73.080 103.165 73.830 103.335 ;
        RECT 73.075 102.615 73.405 102.995 ;
        RECT 73.575 102.875 73.830 103.165 ;
        RECT 74.005 102.615 75.675 103.385 ;
        RECT 76.360 103.435 76.770 103.985 ;
        RECT 78.640 103.825 78.810 104.445 ;
        RECT 80.030 104.275 80.200 104.655 ;
        RECT 81.135 104.535 81.305 104.995 ;
        RECT 81.475 104.705 81.845 105.165 ;
        RECT 82.140 104.565 82.310 104.905 ;
        RECT 82.480 104.735 82.810 105.165 ;
        RECT 83.045 104.565 83.215 104.905 ;
        RECT 78.980 104.105 80.200 104.275 ;
        RECT 80.370 104.195 80.830 104.485 ;
        RECT 81.135 104.365 81.695 104.535 ;
        RECT 82.140 104.395 83.215 104.565 ;
        RECT 83.385 104.665 84.065 104.995 ;
        RECT 84.280 104.665 84.530 104.995 ;
        RECT 84.700 104.705 84.950 105.165 ;
        RECT 81.525 104.225 81.695 104.365 ;
        RECT 80.370 104.185 81.335 104.195 ;
        RECT 80.030 104.015 80.200 104.105 ;
        RECT 80.660 104.025 81.335 104.185 ;
        RECT 78.640 103.815 78.985 103.825 ;
        RECT 76.955 103.605 78.985 103.815 ;
        RECT 75.845 102.615 76.135 103.340 ;
        RECT 76.360 103.265 78.125 103.435 ;
        RECT 76.615 102.615 76.785 103.085 ;
        RECT 76.955 102.785 77.285 103.265 ;
        RECT 77.455 102.615 77.625 103.085 ;
        RECT 77.795 102.785 78.125 103.265 ;
        RECT 78.295 102.615 78.465 103.425 ;
        RECT 78.660 103.350 78.985 103.605 ;
        RECT 78.665 102.995 78.985 103.350 ;
        RECT 79.155 103.565 79.695 103.935 ;
        RECT 80.030 103.845 80.435 104.015 ;
        RECT 79.155 103.165 79.395 103.565 ;
        RECT 79.875 103.395 80.095 103.675 ;
        RECT 79.565 103.225 80.095 103.395 ;
        RECT 79.565 102.995 79.735 103.225 ;
        RECT 80.265 103.065 80.435 103.845 ;
        RECT 80.605 103.235 80.955 103.855 ;
        RECT 81.125 103.235 81.335 104.025 ;
        RECT 81.525 104.055 83.025 104.225 ;
        RECT 81.525 103.365 81.695 104.055 ;
        RECT 83.385 103.885 83.555 104.665 ;
        RECT 84.360 104.535 84.530 104.665 ;
        RECT 81.865 103.715 83.555 103.885 ;
        RECT 83.725 104.105 84.190 104.495 ;
        RECT 84.360 104.365 84.755 104.535 ;
        RECT 81.865 103.535 82.035 103.715 ;
        RECT 78.665 102.825 79.735 102.995 ;
        RECT 79.905 102.615 80.095 103.055 ;
        RECT 80.265 102.785 81.215 103.065 ;
        RECT 81.525 102.975 81.785 103.365 ;
        RECT 82.205 103.295 82.995 103.545 ;
        RECT 81.435 102.805 81.785 102.975 ;
        RECT 81.995 102.615 82.325 103.075 ;
        RECT 83.200 103.005 83.370 103.715 ;
        RECT 83.725 103.515 83.895 104.105 ;
        RECT 83.540 103.295 83.895 103.515 ;
        RECT 84.065 103.295 84.415 103.915 ;
        RECT 84.585 103.005 84.755 104.365 ;
        RECT 85.120 104.195 85.445 104.980 ;
        RECT 84.925 103.145 85.385 104.195 ;
        RECT 83.200 102.835 84.055 103.005 ;
        RECT 84.260 102.835 84.755 103.005 ;
        RECT 84.925 102.615 85.255 102.975 ;
        RECT 85.615 102.875 85.785 104.995 ;
        RECT 85.955 104.665 86.285 105.165 ;
        RECT 86.455 104.495 86.710 104.995 ;
        RECT 85.960 104.325 86.710 104.495 ;
        RECT 87.195 104.325 87.365 105.165 ;
        RECT 85.960 103.335 86.190 104.325 ;
        RECT 87.575 104.155 87.825 104.995 ;
        RECT 88.035 104.325 88.205 105.165 ;
        RECT 88.375 104.155 88.665 104.995 ;
        RECT 86.360 103.505 86.710 104.155 ;
        RECT 86.940 103.985 88.665 104.155 ;
        RECT 88.875 104.105 89.045 105.165 ;
        RECT 89.340 104.785 89.670 105.165 ;
        RECT 89.850 104.615 90.020 104.905 ;
        RECT 90.190 104.705 90.440 105.165 ;
        RECT 89.220 104.445 90.020 104.615 ;
        RECT 90.610 104.655 91.480 104.995 ;
        RECT 86.940 103.435 87.350 103.985 ;
        RECT 89.220 103.825 89.390 104.445 ;
        RECT 90.610 104.275 90.780 104.655 ;
        RECT 91.715 104.535 91.885 104.995 ;
        RECT 92.055 104.705 92.425 105.165 ;
        RECT 92.720 104.565 92.890 104.905 ;
        RECT 93.060 104.735 93.390 105.165 ;
        RECT 93.625 104.565 93.795 104.905 ;
        RECT 89.560 104.105 90.780 104.275 ;
        RECT 90.950 104.195 91.410 104.485 ;
        RECT 91.715 104.365 92.275 104.535 ;
        RECT 92.720 104.395 93.795 104.565 ;
        RECT 93.965 104.665 94.645 104.995 ;
        RECT 94.860 104.665 95.110 104.995 ;
        RECT 95.280 104.705 95.530 105.165 ;
        RECT 92.105 104.225 92.275 104.365 ;
        RECT 90.950 104.185 91.915 104.195 ;
        RECT 90.610 104.015 90.780 104.105 ;
        RECT 91.240 104.025 91.915 104.185 ;
        RECT 89.220 103.815 89.565 103.825 ;
        RECT 87.535 103.605 89.565 103.815 ;
        RECT 85.960 103.165 86.710 103.335 ;
        RECT 86.940 103.265 88.705 103.435 ;
        RECT 85.955 102.615 86.285 102.995 ;
        RECT 86.455 102.875 86.710 103.165 ;
        RECT 87.195 102.615 87.365 103.085 ;
        RECT 87.535 102.785 87.865 103.265 ;
        RECT 88.035 102.615 88.205 103.085 ;
        RECT 88.375 102.785 88.705 103.265 ;
        RECT 88.875 102.615 89.045 103.425 ;
        RECT 89.240 103.350 89.565 103.605 ;
        RECT 89.245 102.995 89.565 103.350 ;
        RECT 89.735 103.565 90.275 103.935 ;
        RECT 90.610 103.845 91.015 104.015 ;
        RECT 89.735 103.165 89.975 103.565 ;
        RECT 90.455 103.395 90.675 103.675 ;
        RECT 90.145 103.225 90.675 103.395 ;
        RECT 90.145 102.995 90.315 103.225 ;
        RECT 90.845 103.065 91.015 103.845 ;
        RECT 91.185 103.235 91.535 103.855 ;
        RECT 91.705 103.235 91.915 104.025 ;
        RECT 92.105 104.055 93.605 104.225 ;
        RECT 92.105 103.365 92.275 104.055 ;
        RECT 93.965 103.885 94.135 104.665 ;
        RECT 94.940 104.535 95.110 104.665 ;
        RECT 92.445 103.715 94.135 103.885 ;
        RECT 94.305 104.105 94.770 104.495 ;
        RECT 94.940 104.365 95.335 104.535 ;
        RECT 92.445 103.535 92.615 103.715 ;
        RECT 89.245 102.825 90.315 102.995 ;
        RECT 90.485 102.615 90.675 103.055 ;
        RECT 90.845 102.785 91.795 103.065 ;
        RECT 92.105 102.975 92.365 103.365 ;
        RECT 92.785 103.295 93.575 103.545 ;
        RECT 92.015 102.805 92.365 102.975 ;
        RECT 92.575 102.615 92.905 103.075 ;
        RECT 93.780 103.005 93.950 103.715 ;
        RECT 94.305 103.515 94.475 104.105 ;
        RECT 94.120 103.295 94.475 103.515 ;
        RECT 94.645 103.295 94.995 103.915 ;
        RECT 95.165 103.005 95.335 104.365 ;
        RECT 95.700 104.195 96.025 104.980 ;
        RECT 95.505 103.145 95.965 104.195 ;
        RECT 93.780 102.835 94.635 103.005 ;
        RECT 94.840 102.835 95.335 103.005 ;
        RECT 95.505 102.615 95.835 102.975 ;
        RECT 96.195 102.875 96.365 104.995 ;
        RECT 96.535 104.665 96.865 105.165 ;
        RECT 97.035 104.495 97.290 104.995 ;
        RECT 96.540 104.325 97.290 104.495 ;
        RECT 96.540 103.335 96.770 104.325 ;
        RECT 96.940 103.505 97.290 104.155 ;
        RECT 97.925 104.075 101.435 105.165 ;
        RECT 97.925 103.555 99.615 104.075 ;
        RECT 101.605 104.000 101.895 105.165 ;
        RECT 102.375 104.325 102.545 105.165 ;
        RECT 102.755 104.155 103.005 104.995 ;
        RECT 103.215 104.325 103.385 105.165 ;
        RECT 103.555 104.155 103.845 104.995 ;
        RECT 102.120 103.985 103.845 104.155 ;
        RECT 104.055 104.105 104.225 105.165 ;
        RECT 104.520 104.785 104.850 105.165 ;
        RECT 105.030 104.615 105.200 104.905 ;
        RECT 105.370 104.705 105.620 105.165 ;
        RECT 104.400 104.445 105.200 104.615 ;
        RECT 105.790 104.655 106.660 104.995 ;
        RECT 99.785 103.385 101.435 103.905 ;
        RECT 96.540 103.165 97.290 103.335 ;
        RECT 96.535 102.615 96.865 102.995 ;
        RECT 97.035 102.875 97.290 103.165 ;
        RECT 97.925 102.615 101.435 103.385 ;
        RECT 102.120 103.435 102.530 103.985 ;
        RECT 104.400 103.825 104.570 104.445 ;
        RECT 105.790 104.275 105.960 104.655 ;
        RECT 106.895 104.535 107.065 104.995 ;
        RECT 107.235 104.705 107.605 105.165 ;
        RECT 107.900 104.565 108.070 104.905 ;
        RECT 108.240 104.735 108.570 105.165 ;
        RECT 108.805 104.565 108.975 104.905 ;
        RECT 104.740 104.105 105.960 104.275 ;
        RECT 106.130 104.195 106.590 104.485 ;
        RECT 106.895 104.365 107.455 104.535 ;
        RECT 107.900 104.395 108.975 104.565 ;
        RECT 109.145 104.665 109.825 104.995 ;
        RECT 110.040 104.665 110.290 104.995 ;
        RECT 110.460 104.705 110.710 105.165 ;
        RECT 107.285 104.225 107.455 104.365 ;
        RECT 106.130 104.185 107.095 104.195 ;
        RECT 105.790 104.015 105.960 104.105 ;
        RECT 106.420 104.025 107.095 104.185 ;
        RECT 104.400 103.815 104.745 103.825 ;
        RECT 102.715 103.605 104.745 103.815 ;
        RECT 101.605 102.615 101.895 103.340 ;
        RECT 102.120 103.265 103.885 103.435 ;
        RECT 102.375 102.615 102.545 103.085 ;
        RECT 102.715 102.785 103.045 103.265 ;
        RECT 103.215 102.615 103.385 103.085 ;
        RECT 103.555 102.785 103.885 103.265 ;
        RECT 104.055 102.615 104.225 103.425 ;
        RECT 104.420 103.350 104.745 103.605 ;
        RECT 104.425 102.995 104.745 103.350 ;
        RECT 104.915 103.565 105.455 103.935 ;
        RECT 105.790 103.845 106.195 104.015 ;
        RECT 104.915 103.165 105.155 103.565 ;
        RECT 105.635 103.395 105.855 103.675 ;
        RECT 105.325 103.225 105.855 103.395 ;
        RECT 105.325 102.995 105.495 103.225 ;
        RECT 106.025 103.065 106.195 103.845 ;
        RECT 106.365 103.235 106.715 103.855 ;
        RECT 106.885 103.235 107.095 104.025 ;
        RECT 107.285 104.055 108.785 104.225 ;
        RECT 107.285 103.365 107.455 104.055 ;
        RECT 109.145 103.885 109.315 104.665 ;
        RECT 110.120 104.535 110.290 104.665 ;
        RECT 107.625 103.715 109.315 103.885 ;
        RECT 109.485 104.105 109.950 104.495 ;
        RECT 110.120 104.365 110.515 104.535 ;
        RECT 107.625 103.535 107.795 103.715 ;
        RECT 104.425 102.825 105.495 102.995 ;
        RECT 105.665 102.615 105.855 103.055 ;
        RECT 106.025 102.785 106.975 103.065 ;
        RECT 107.285 102.975 107.545 103.365 ;
        RECT 107.965 103.295 108.755 103.545 ;
        RECT 107.195 102.805 107.545 102.975 ;
        RECT 107.755 102.615 108.085 103.075 ;
        RECT 108.960 103.005 109.130 103.715 ;
        RECT 109.485 103.515 109.655 104.105 ;
        RECT 109.300 103.295 109.655 103.515 ;
        RECT 109.825 103.295 110.175 103.915 ;
        RECT 110.345 103.005 110.515 104.365 ;
        RECT 110.880 104.195 111.205 104.980 ;
        RECT 110.685 103.145 111.145 104.195 ;
        RECT 108.960 102.835 109.815 103.005 ;
        RECT 110.020 102.835 110.515 103.005 ;
        RECT 110.685 102.615 111.015 102.975 ;
        RECT 111.375 102.875 111.545 104.995 ;
        RECT 111.715 104.665 112.045 105.165 ;
        RECT 112.215 104.495 112.470 104.995 ;
        RECT 111.720 104.325 112.470 104.495 ;
        RECT 112.650 104.495 112.905 104.995 ;
        RECT 113.075 104.665 113.405 105.165 ;
        RECT 112.650 104.325 113.400 104.495 ;
        RECT 111.720 103.335 111.950 104.325 ;
        RECT 112.120 103.505 112.470 104.155 ;
        RECT 112.650 103.505 113.000 104.155 ;
        RECT 113.170 103.335 113.400 104.325 ;
        RECT 111.720 103.165 112.470 103.335 ;
        RECT 111.715 102.615 112.045 102.995 ;
        RECT 112.215 102.875 112.470 103.165 ;
        RECT 112.650 103.165 113.400 103.335 ;
        RECT 112.650 102.875 112.905 103.165 ;
        RECT 113.075 102.615 113.405 102.995 ;
        RECT 113.575 102.875 113.745 104.995 ;
        RECT 113.915 104.195 114.240 104.980 ;
        RECT 114.410 104.705 114.660 105.165 ;
        RECT 114.830 104.665 115.080 104.995 ;
        RECT 115.295 104.665 115.975 104.995 ;
        RECT 114.830 104.535 115.000 104.665 ;
        RECT 114.605 104.365 115.000 104.535 ;
        RECT 113.975 103.145 114.435 104.195 ;
        RECT 114.605 103.005 114.775 104.365 ;
        RECT 115.170 104.105 115.635 104.495 ;
        RECT 114.945 103.295 115.295 103.915 ;
        RECT 115.465 103.515 115.635 104.105 ;
        RECT 115.805 103.885 115.975 104.665 ;
        RECT 116.145 104.565 116.315 104.905 ;
        RECT 116.550 104.735 116.880 105.165 ;
        RECT 117.050 104.565 117.220 104.905 ;
        RECT 117.515 104.705 117.885 105.165 ;
        RECT 116.145 104.395 117.220 104.565 ;
        RECT 118.055 104.535 118.225 104.995 ;
        RECT 118.460 104.655 119.330 104.995 ;
        RECT 119.500 104.705 119.750 105.165 ;
        RECT 117.665 104.365 118.225 104.535 ;
        RECT 117.665 104.225 117.835 104.365 ;
        RECT 116.335 104.055 117.835 104.225 ;
        RECT 118.530 104.195 118.990 104.485 ;
        RECT 115.805 103.715 117.495 103.885 ;
        RECT 115.465 103.295 115.820 103.515 ;
        RECT 115.990 103.005 116.160 103.715 ;
        RECT 116.365 103.295 117.155 103.545 ;
        RECT 117.325 103.535 117.495 103.715 ;
        RECT 117.665 103.365 117.835 104.055 ;
        RECT 114.105 102.615 114.435 102.975 ;
        RECT 114.605 102.835 115.100 103.005 ;
        RECT 115.305 102.835 116.160 103.005 ;
        RECT 117.035 102.615 117.365 103.075 ;
        RECT 117.575 102.975 117.835 103.365 ;
        RECT 118.025 104.185 118.990 104.195 ;
        RECT 119.160 104.275 119.330 104.655 ;
        RECT 119.920 104.615 120.090 104.905 ;
        RECT 120.270 104.785 120.600 105.165 ;
        RECT 119.920 104.445 120.720 104.615 ;
        RECT 118.025 104.025 118.700 104.185 ;
        RECT 119.160 104.105 120.380 104.275 ;
        RECT 118.025 103.235 118.235 104.025 ;
        RECT 119.160 104.015 119.330 104.105 ;
        RECT 118.405 103.235 118.755 103.855 ;
        RECT 118.925 103.845 119.330 104.015 ;
        RECT 118.925 103.065 119.095 103.845 ;
        RECT 119.265 103.395 119.485 103.675 ;
        RECT 119.665 103.565 120.205 103.935 ;
        RECT 120.550 103.825 120.720 104.445 ;
        RECT 120.895 104.105 121.065 105.165 ;
        RECT 121.275 104.155 121.565 104.995 ;
        RECT 121.735 104.325 121.905 105.165 ;
        RECT 122.115 104.155 122.365 104.995 ;
        RECT 122.575 104.325 122.745 105.165 ;
        RECT 121.275 103.985 123.000 104.155 ;
        RECT 119.265 103.225 119.795 103.395 ;
        RECT 117.575 102.805 117.925 102.975 ;
        RECT 118.145 102.785 119.095 103.065 ;
        RECT 119.265 102.615 119.455 103.055 ;
        RECT 119.625 102.995 119.795 103.225 ;
        RECT 119.965 103.165 120.205 103.565 ;
        RECT 120.375 103.815 120.720 103.825 ;
        RECT 120.375 103.605 122.405 103.815 ;
        RECT 120.375 103.350 120.700 103.605 ;
        RECT 122.590 103.435 123.000 103.985 ;
        RECT 123.225 104.075 124.895 105.165 ;
        RECT 125.065 104.090 125.335 104.995 ;
        RECT 125.505 104.405 125.835 105.165 ;
        RECT 126.015 104.235 126.195 104.995 ;
        RECT 123.225 103.555 123.975 104.075 ;
        RECT 120.375 102.995 120.695 103.350 ;
        RECT 119.625 102.825 120.695 102.995 ;
        RECT 120.895 102.615 121.065 103.425 ;
        RECT 121.235 103.265 123.000 103.435 ;
        RECT 124.145 103.385 124.895 103.905 ;
        RECT 121.235 102.785 121.565 103.265 ;
        RECT 121.735 102.615 121.905 103.085 ;
        RECT 122.075 102.785 122.405 103.265 ;
        RECT 122.575 102.615 122.745 103.085 ;
        RECT 123.225 102.615 124.895 103.385 ;
        RECT 125.065 103.290 125.245 104.090 ;
        RECT 125.520 104.065 126.195 104.235 ;
        RECT 126.445 104.075 127.655 105.165 ;
        RECT 125.520 103.920 125.690 104.065 ;
        RECT 125.415 103.590 125.690 103.920 ;
        RECT 125.520 103.335 125.690 103.590 ;
        RECT 125.915 103.515 126.255 103.885 ;
        RECT 126.445 103.535 126.965 104.075 ;
        RECT 127.135 103.365 127.655 103.905 ;
        RECT 125.065 102.785 125.325 103.290 ;
        RECT 125.520 103.165 126.185 103.335 ;
        RECT 125.505 102.615 125.835 102.995 ;
        RECT 126.015 102.785 126.185 103.165 ;
        RECT 126.445 102.615 127.655 103.365 ;
        RECT 14.580 102.445 127.740 102.615 ;
        RECT 14.665 101.695 15.875 102.445 ;
        RECT 14.665 101.155 15.185 101.695 ;
        RECT 16.045 101.675 18.635 102.445 ;
        RECT 18.810 101.900 24.155 102.445 ;
        RECT 15.355 100.985 15.875 101.525 ;
        RECT 14.665 99.895 15.875 100.985 ;
        RECT 16.045 100.985 17.255 101.505 ;
        RECT 17.425 101.155 18.635 101.675 ;
        RECT 16.045 99.895 18.635 100.985 ;
        RECT 20.400 100.330 20.750 101.580 ;
        RECT 22.230 101.070 22.570 101.900 ;
        RECT 24.325 101.720 24.615 102.445 ;
        RECT 25.095 101.975 25.265 102.445 ;
        RECT 25.435 101.795 25.765 102.275 ;
        RECT 25.935 101.975 26.105 102.445 ;
        RECT 26.275 101.795 26.605 102.275 ;
        RECT 24.840 101.625 26.605 101.795 ;
        RECT 26.775 101.635 26.945 102.445 ;
        RECT 27.145 102.065 28.215 102.235 ;
        RECT 27.145 101.710 27.465 102.065 ;
        RECT 24.840 101.075 25.250 101.625 ;
        RECT 27.140 101.455 27.465 101.710 ;
        RECT 25.435 101.245 27.465 101.455 ;
        RECT 27.120 101.235 27.465 101.245 ;
        RECT 27.635 101.495 27.875 101.895 ;
        RECT 28.045 101.835 28.215 102.065 ;
        RECT 28.385 102.005 28.575 102.445 ;
        RECT 28.745 101.995 29.695 102.275 ;
        RECT 29.915 102.085 30.265 102.255 ;
        RECT 28.045 101.665 28.575 101.835 ;
        RECT 18.810 99.895 24.155 100.330 ;
        RECT 24.325 99.895 24.615 101.060 ;
        RECT 24.840 100.905 26.565 101.075 ;
        RECT 25.095 99.895 25.265 100.735 ;
        RECT 25.475 100.065 25.725 100.905 ;
        RECT 25.935 99.895 26.105 100.735 ;
        RECT 26.275 100.065 26.565 100.905 ;
        RECT 26.775 99.895 26.945 100.955 ;
        RECT 27.120 100.615 27.290 101.235 ;
        RECT 27.635 101.125 28.175 101.495 ;
        RECT 28.355 101.385 28.575 101.665 ;
        RECT 28.745 101.215 28.915 101.995 ;
        RECT 28.510 101.045 28.915 101.215 ;
        RECT 29.085 101.205 29.435 101.825 ;
        RECT 28.510 100.955 28.680 101.045 ;
        RECT 29.605 101.035 29.815 101.825 ;
        RECT 27.460 100.785 28.680 100.955 ;
        RECT 29.140 100.875 29.815 101.035 ;
        RECT 27.120 100.445 27.920 100.615 ;
        RECT 27.240 99.895 27.570 100.275 ;
        RECT 27.750 100.155 27.920 100.445 ;
        RECT 28.510 100.405 28.680 100.785 ;
        RECT 28.850 100.865 29.815 100.875 ;
        RECT 30.005 101.695 30.265 102.085 ;
        RECT 30.475 101.985 30.805 102.445 ;
        RECT 31.680 102.055 32.535 102.225 ;
        RECT 32.740 102.055 33.235 102.225 ;
        RECT 33.405 102.085 33.735 102.445 ;
        RECT 30.005 101.005 30.175 101.695 ;
        RECT 30.345 101.345 30.515 101.525 ;
        RECT 30.685 101.515 31.475 101.765 ;
        RECT 31.680 101.345 31.850 102.055 ;
        RECT 32.020 101.545 32.375 101.765 ;
        RECT 30.345 101.175 32.035 101.345 ;
        RECT 28.850 100.575 29.310 100.865 ;
        RECT 30.005 100.835 31.505 101.005 ;
        RECT 30.005 100.695 30.175 100.835 ;
        RECT 29.615 100.525 30.175 100.695 ;
        RECT 28.090 99.895 28.340 100.355 ;
        RECT 28.510 100.065 29.380 100.405 ;
        RECT 29.615 100.065 29.785 100.525 ;
        RECT 30.620 100.495 31.695 100.665 ;
        RECT 29.955 99.895 30.325 100.355 ;
        RECT 30.620 100.155 30.790 100.495 ;
        RECT 30.960 99.895 31.290 100.325 ;
        RECT 31.525 100.155 31.695 100.495 ;
        RECT 31.865 100.395 32.035 101.175 ;
        RECT 32.205 100.955 32.375 101.545 ;
        RECT 32.545 101.145 32.895 101.765 ;
        RECT 32.205 100.565 32.670 100.955 ;
        RECT 33.065 100.695 33.235 102.055 ;
        RECT 33.405 100.865 33.865 101.915 ;
        RECT 32.840 100.525 33.235 100.695 ;
        RECT 32.840 100.395 33.010 100.525 ;
        RECT 31.865 100.065 32.545 100.395 ;
        RECT 32.760 100.065 33.010 100.395 ;
        RECT 33.180 99.895 33.430 100.355 ;
        RECT 33.600 100.080 33.925 100.865 ;
        RECT 34.095 100.065 34.265 102.185 ;
        RECT 34.435 102.065 34.765 102.445 ;
        RECT 34.935 101.895 35.190 102.185 ;
        RECT 34.440 101.725 35.190 101.895 ;
        RECT 34.440 100.735 34.670 101.725 ;
        RECT 35.365 101.675 37.035 102.445 ;
        RECT 37.205 101.720 37.495 102.445 ;
        RECT 37.665 101.695 38.875 102.445 ;
        RECT 39.050 101.900 44.395 102.445 ;
        RECT 44.570 101.900 49.915 102.445 ;
        RECT 34.840 100.905 35.190 101.555 ;
        RECT 35.365 100.985 36.115 101.505 ;
        RECT 36.285 101.155 37.035 101.675 ;
        RECT 34.440 100.565 35.190 100.735 ;
        RECT 34.435 99.895 34.765 100.395 ;
        RECT 34.935 100.065 35.190 100.565 ;
        RECT 35.365 99.895 37.035 100.985 ;
        RECT 37.205 99.895 37.495 101.060 ;
        RECT 37.665 100.985 38.185 101.525 ;
        RECT 38.355 101.155 38.875 101.695 ;
        RECT 37.665 99.895 38.875 100.985 ;
        RECT 40.640 100.330 40.990 101.580 ;
        RECT 42.470 101.070 42.810 101.900 ;
        RECT 46.160 100.330 46.510 101.580 ;
        RECT 47.990 101.070 48.330 101.900 ;
        RECT 50.085 101.720 50.375 102.445 ;
        RECT 50.545 101.695 51.755 102.445 ;
        RECT 51.930 101.900 57.275 102.445 ;
        RECT 57.450 101.900 62.795 102.445 ;
        RECT 39.050 99.895 44.395 100.330 ;
        RECT 44.570 99.895 49.915 100.330 ;
        RECT 50.085 99.895 50.375 101.060 ;
        RECT 50.545 100.985 51.065 101.525 ;
        RECT 51.235 101.155 51.755 101.695 ;
        RECT 50.545 99.895 51.755 100.985 ;
        RECT 53.520 100.330 53.870 101.580 ;
        RECT 55.350 101.070 55.690 101.900 ;
        RECT 59.040 100.330 59.390 101.580 ;
        RECT 60.870 101.070 61.210 101.900 ;
        RECT 62.965 101.720 63.255 102.445 ;
        RECT 63.425 101.695 64.635 102.445 ;
        RECT 64.810 101.900 70.155 102.445 ;
        RECT 70.330 101.900 75.675 102.445 ;
        RECT 51.930 99.895 57.275 100.330 ;
        RECT 57.450 99.895 62.795 100.330 ;
        RECT 62.965 99.895 63.255 101.060 ;
        RECT 63.425 100.985 63.945 101.525 ;
        RECT 64.115 101.155 64.635 101.695 ;
        RECT 63.425 99.895 64.635 100.985 ;
        RECT 66.400 100.330 66.750 101.580 ;
        RECT 68.230 101.070 68.570 101.900 ;
        RECT 71.920 100.330 72.270 101.580 ;
        RECT 73.750 101.070 74.090 101.900 ;
        RECT 75.845 101.720 76.135 102.445 ;
        RECT 76.305 101.695 77.515 102.445 ;
        RECT 77.690 101.900 83.035 102.445 ;
        RECT 83.210 101.900 88.555 102.445 ;
        RECT 64.810 99.895 70.155 100.330 ;
        RECT 70.330 99.895 75.675 100.330 ;
        RECT 75.845 99.895 76.135 101.060 ;
        RECT 76.305 100.985 76.825 101.525 ;
        RECT 76.995 101.155 77.515 101.695 ;
        RECT 76.305 99.895 77.515 100.985 ;
        RECT 79.280 100.330 79.630 101.580 ;
        RECT 81.110 101.070 81.450 101.900 ;
        RECT 84.800 100.330 85.150 101.580 ;
        RECT 86.630 101.070 86.970 101.900 ;
        RECT 88.725 101.720 89.015 102.445 ;
        RECT 89.185 101.675 90.855 102.445 ;
        RECT 91.335 101.975 91.505 102.445 ;
        RECT 91.675 101.795 92.005 102.275 ;
        RECT 92.175 101.975 92.345 102.445 ;
        RECT 92.515 101.795 92.845 102.275 ;
        RECT 77.690 99.895 83.035 100.330 ;
        RECT 83.210 99.895 88.555 100.330 ;
        RECT 88.725 99.895 89.015 101.060 ;
        RECT 89.185 100.985 89.935 101.505 ;
        RECT 90.105 101.155 90.855 101.675 ;
        RECT 91.080 101.625 92.845 101.795 ;
        RECT 93.015 101.635 93.185 102.445 ;
        RECT 93.385 102.065 94.455 102.235 ;
        RECT 93.385 101.710 93.705 102.065 ;
        RECT 91.080 101.075 91.490 101.625 ;
        RECT 93.380 101.455 93.705 101.710 ;
        RECT 91.675 101.245 93.705 101.455 ;
        RECT 93.360 101.235 93.705 101.245 ;
        RECT 93.875 101.495 94.115 101.895 ;
        RECT 94.285 101.835 94.455 102.065 ;
        RECT 94.625 102.005 94.815 102.445 ;
        RECT 94.985 101.995 95.935 102.275 ;
        RECT 96.155 102.085 96.505 102.255 ;
        RECT 94.285 101.665 94.815 101.835 ;
        RECT 89.185 99.895 90.855 100.985 ;
        RECT 91.080 100.905 92.805 101.075 ;
        RECT 91.335 99.895 91.505 100.735 ;
        RECT 91.715 100.065 91.965 100.905 ;
        RECT 92.175 99.895 92.345 100.735 ;
        RECT 92.515 100.065 92.805 100.905 ;
        RECT 93.015 99.895 93.185 100.955 ;
        RECT 93.360 100.615 93.530 101.235 ;
        RECT 93.875 101.125 94.415 101.495 ;
        RECT 94.595 101.385 94.815 101.665 ;
        RECT 94.985 101.215 95.155 101.995 ;
        RECT 94.750 101.045 95.155 101.215 ;
        RECT 95.325 101.205 95.675 101.825 ;
        RECT 94.750 100.955 94.920 101.045 ;
        RECT 95.845 101.035 96.055 101.825 ;
        RECT 93.700 100.785 94.920 100.955 ;
        RECT 95.380 100.875 96.055 101.035 ;
        RECT 93.360 100.445 94.160 100.615 ;
        RECT 93.480 99.895 93.810 100.275 ;
        RECT 93.990 100.155 94.160 100.445 ;
        RECT 94.750 100.405 94.920 100.785 ;
        RECT 95.090 100.865 96.055 100.875 ;
        RECT 96.245 101.695 96.505 102.085 ;
        RECT 96.715 101.985 97.045 102.445 ;
        RECT 97.920 102.055 98.775 102.225 ;
        RECT 98.980 102.055 99.475 102.225 ;
        RECT 99.645 102.085 99.975 102.445 ;
        RECT 96.245 101.005 96.415 101.695 ;
        RECT 96.585 101.345 96.755 101.525 ;
        RECT 96.925 101.515 97.715 101.765 ;
        RECT 97.920 101.345 98.090 102.055 ;
        RECT 98.260 101.545 98.615 101.765 ;
        RECT 96.585 101.175 98.275 101.345 ;
        RECT 95.090 100.575 95.550 100.865 ;
        RECT 96.245 100.835 97.745 101.005 ;
        RECT 96.245 100.695 96.415 100.835 ;
        RECT 95.855 100.525 96.415 100.695 ;
        RECT 94.330 99.895 94.580 100.355 ;
        RECT 94.750 100.065 95.620 100.405 ;
        RECT 95.855 100.065 96.025 100.525 ;
        RECT 96.860 100.495 97.935 100.665 ;
        RECT 96.195 99.895 96.565 100.355 ;
        RECT 96.860 100.155 97.030 100.495 ;
        RECT 97.200 99.895 97.530 100.325 ;
        RECT 97.765 100.155 97.935 100.495 ;
        RECT 98.105 100.395 98.275 101.175 ;
        RECT 98.445 100.955 98.615 101.545 ;
        RECT 98.785 101.145 99.135 101.765 ;
        RECT 98.445 100.565 98.910 100.955 ;
        RECT 99.305 100.695 99.475 102.055 ;
        RECT 99.645 100.865 100.105 101.915 ;
        RECT 99.080 100.525 99.475 100.695 ;
        RECT 99.080 100.395 99.250 100.525 ;
        RECT 98.105 100.065 98.785 100.395 ;
        RECT 99.000 100.065 99.250 100.395 ;
        RECT 99.420 99.895 99.670 100.355 ;
        RECT 99.840 100.080 100.165 100.865 ;
        RECT 100.335 100.065 100.505 102.185 ;
        RECT 100.675 102.065 101.005 102.445 ;
        RECT 101.175 101.895 101.430 102.185 ;
        RECT 100.680 101.725 101.430 101.895 ;
        RECT 100.680 100.735 100.910 101.725 ;
        RECT 101.605 101.720 101.895 102.445 ;
        RECT 102.065 101.695 103.275 102.445 ;
        RECT 103.450 101.900 108.795 102.445 ;
        RECT 108.970 101.900 114.315 102.445 ;
        RECT 101.080 100.905 101.430 101.555 ;
        RECT 100.680 100.565 101.430 100.735 ;
        RECT 100.675 99.895 101.005 100.395 ;
        RECT 101.175 100.065 101.430 100.565 ;
        RECT 101.605 99.895 101.895 101.060 ;
        RECT 102.065 100.985 102.585 101.525 ;
        RECT 102.755 101.155 103.275 101.695 ;
        RECT 102.065 99.895 103.275 100.985 ;
        RECT 105.040 100.330 105.390 101.580 ;
        RECT 106.870 101.070 107.210 101.900 ;
        RECT 110.560 100.330 110.910 101.580 ;
        RECT 112.390 101.070 112.730 101.900 ;
        RECT 114.485 101.720 114.775 102.445 ;
        RECT 115.865 101.675 119.375 102.445 ;
        RECT 103.450 99.895 108.795 100.330 ;
        RECT 108.970 99.895 114.315 100.330 ;
        RECT 114.485 99.895 114.775 101.060 ;
        RECT 115.865 100.985 117.555 101.505 ;
        RECT 117.725 101.155 119.375 101.675 ;
        RECT 119.585 101.625 119.815 102.445 ;
        RECT 119.985 101.645 120.315 102.275 ;
        RECT 119.565 101.205 119.895 101.455 ;
        RECT 120.065 101.045 120.315 101.645 ;
        RECT 120.485 101.625 120.695 102.445 ;
        RECT 120.930 101.900 126.275 102.445 ;
        RECT 115.865 99.895 119.375 100.985 ;
        RECT 119.585 99.895 119.815 101.035 ;
        RECT 119.985 100.065 120.315 101.045 ;
        RECT 120.485 99.895 120.695 101.035 ;
        RECT 122.520 100.330 122.870 101.580 ;
        RECT 124.350 101.070 124.690 101.900 ;
        RECT 126.445 101.695 127.655 102.445 ;
        RECT 126.445 100.985 126.965 101.525 ;
        RECT 127.135 101.155 127.655 101.695 ;
        RECT 120.930 99.895 126.275 100.330 ;
        RECT 126.445 99.895 127.655 100.985 ;
        RECT 14.580 99.725 127.740 99.895 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.580 211.090 127.740 211.570 ;
        RECT 14.580 208.370 127.740 208.850 ;
        RECT 73.530 207.830 73.850 207.890 ;
        RECT 74.925 207.830 75.215 207.875 ;
        RECT 73.530 207.690 79.280 207.830 ;
        RECT 73.530 207.630 73.850 207.690 ;
        RECT 74.925 207.645 75.215 207.690 ;
        RECT 66.170 207.150 66.490 207.210 ;
        RECT 72.625 207.150 72.915 207.195 ;
        RECT 66.170 207.010 72.915 207.150 ;
        RECT 66.170 206.950 66.490 207.010 ;
        RECT 72.625 206.965 72.915 207.010 ;
        RECT 73.070 207.150 73.390 207.210 ;
        RECT 79.140 207.195 79.280 207.690 ;
        RECT 79.510 207.290 79.830 207.550 ;
        RECT 74.005 207.150 74.295 207.195 ;
        RECT 73.070 207.010 74.295 207.150 ;
        RECT 73.070 206.950 73.390 207.010 ;
        RECT 74.005 206.965 74.295 207.010 ;
        RECT 79.065 206.965 79.355 207.195 ;
        RECT 73.085 206.470 73.375 206.515 ;
        RECT 73.990 206.470 74.310 206.530 ;
        RECT 73.085 206.330 74.310 206.470 ;
        RECT 73.085 206.285 73.375 206.330 ;
        RECT 73.990 206.270 74.310 206.330 ;
        RECT 75.830 206.470 76.150 206.530 ;
        RECT 77.225 206.470 77.515 206.515 ;
        RECT 75.830 206.330 77.515 206.470 ;
        RECT 75.830 206.270 76.150 206.330 ;
        RECT 77.225 206.285 77.515 206.330 ;
        RECT 14.580 205.650 127.740 206.130 ;
        RECT 73.990 205.450 74.310 205.510 ;
        RECT 73.990 205.310 76.520 205.450 ;
        RECT 73.990 205.250 74.310 205.310 ;
        RECT 67.565 205.110 67.855 205.155 ;
        RECT 69.965 205.110 70.255 205.155 ;
        RECT 73.205 205.110 73.855 205.155 ;
        RECT 67.565 204.970 73.855 205.110 ;
        RECT 67.565 204.925 67.855 204.970 ;
        RECT 69.965 204.925 70.555 204.970 ;
        RECT 73.205 204.925 73.855 204.970 ;
        RECT 65.725 204.770 66.015 204.815 ;
        RECT 66.170 204.770 66.490 204.830 ;
        RECT 67.105 204.770 67.395 204.815 ;
        RECT 65.725 204.630 67.395 204.770 ;
        RECT 65.725 204.585 66.015 204.630 ;
        RECT 66.170 204.570 66.490 204.630 ;
        RECT 67.105 204.585 67.395 204.630 ;
        RECT 70.265 204.610 70.555 204.925 ;
        RECT 75.830 204.910 76.150 205.170 ;
        RECT 76.380 205.110 76.520 205.310 ;
        RECT 79.165 205.110 79.455 205.155 ;
        RECT 82.405 205.110 83.055 205.155 ;
        RECT 76.380 204.970 83.055 205.110 ;
        RECT 79.165 204.925 79.755 204.970 ;
        RECT 82.405 204.925 83.055 204.970 ;
        RECT 83.650 205.110 83.970 205.170 ;
        RECT 85.045 205.110 85.335 205.155 ;
        RECT 83.650 204.970 85.335 205.110 ;
        RECT 71.345 204.770 71.635 204.815 ;
        RECT 74.925 204.770 75.215 204.815 ;
        RECT 76.760 204.770 77.050 204.815 ;
        RECT 71.345 204.630 77.050 204.770 ;
        RECT 71.345 204.585 71.635 204.630 ;
        RECT 74.925 204.585 75.215 204.630 ;
        RECT 76.760 204.585 77.050 204.630 ;
        RECT 79.465 204.610 79.755 204.925 ;
        RECT 83.650 204.910 83.970 204.970 ;
        RECT 85.045 204.925 85.335 204.970 ;
        RECT 80.545 204.770 80.835 204.815 ;
        RECT 84.125 204.770 84.415 204.815 ;
        RECT 85.960 204.770 86.250 204.815 ;
        RECT 80.545 204.630 86.250 204.770 ;
        RECT 80.545 204.585 80.835 204.630 ;
        RECT 84.125 204.585 84.415 204.630 ;
        RECT 85.960 204.585 86.250 204.630 ;
        RECT 63.870 204.430 64.190 204.490 ;
        RECT 77.225 204.430 77.515 204.475 ;
        RECT 63.870 204.290 77.515 204.430 ;
        RECT 63.870 204.230 64.190 204.290 ;
        RECT 77.225 204.245 77.515 204.290 ;
        RECT 86.425 204.430 86.715 204.475 ;
        RECT 88.250 204.430 88.570 204.490 ;
        RECT 86.425 204.290 88.570 204.430 ;
        RECT 86.425 204.245 86.715 204.290 ;
        RECT 88.250 204.230 88.570 204.290 ;
        RECT 71.345 204.090 71.635 204.135 ;
        RECT 74.465 204.090 74.755 204.135 ;
        RECT 76.355 204.090 76.645 204.135 ;
        RECT 71.345 203.950 76.645 204.090 ;
        RECT 71.345 203.905 71.635 203.950 ;
        RECT 74.465 203.905 74.755 203.950 ;
        RECT 76.355 203.905 76.645 203.950 ;
        RECT 80.545 204.090 80.835 204.135 ;
        RECT 83.665 204.090 83.955 204.135 ;
        RECT 85.555 204.090 85.845 204.135 ;
        RECT 80.545 203.950 85.845 204.090 ;
        RECT 80.545 203.905 80.835 203.950 ;
        RECT 83.665 203.905 83.955 203.950 ;
        RECT 85.555 203.905 85.845 203.950 ;
        RECT 64.790 203.750 65.110 203.810 ;
        RECT 65.265 203.750 65.555 203.795 ;
        RECT 64.790 203.610 65.555 203.750 ;
        RECT 64.790 203.550 65.110 203.610 ;
        RECT 65.265 203.565 65.555 203.610 ;
        RECT 68.485 203.750 68.775 203.795 ;
        RECT 73.070 203.750 73.390 203.810 ;
        RECT 68.485 203.610 73.390 203.750 ;
        RECT 68.485 203.565 68.775 203.610 ;
        RECT 73.070 203.550 73.390 203.610 ;
        RECT 73.990 203.750 74.310 203.810 ;
        RECT 77.685 203.750 77.975 203.795 ;
        RECT 73.990 203.610 77.975 203.750 ;
        RECT 73.990 203.550 74.310 203.610 ;
        RECT 77.685 203.565 77.975 203.610 ;
        RECT 14.580 202.930 127.740 203.410 ;
        RECT 63.870 202.730 64.190 202.790 ;
        RECT 60.280 202.590 64.190 202.730 ;
        RECT 59.745 202.050 60.035 202.095 ;
        RECT 60.280 202.050 60.420 202.590 ;
        RECT 63.870 202.530 64.190 202.590 ;
        RECT 66.630 202.730 66.950 202.790 ;
        RECT 70.325 202.730 70.615 202.775 ;
        RECT 66.630 202.590 70.615 202.730 ;
        RECT 66.630 202.530 66.950 202.590 ;
        RECT 70.325 202.545 70.615 202.590 ;
        RECT 77.685 202.545 77.975 202.775 ;
        RECT 60.615 202.390 60.905 202.435 ;
        RECT 62.505 202.390 62.795 202.435 ;
        RECT 65.625 202.390 65.915 202.435 ;
        RECT 76.290 202.390 76.610 202.450 ;
        RECT 77.760 202.390 77.900 202.545 ;
        RECT 60.615 202.250 65.915 202.390 ;
        RECT 60.615 202.205 60.905 202.250 ;
        RECT 62.505 202.205 62.795 202.250 ;
        RECT 65.625 202.205 65.915 202.250 ;
        RECT 69.940 202.250 73.760 202.390 ;
        RECT 59.745 201.910 60.420 202.050 ;
        RECT 59.745 201.865 60.035 201.910 ;
        RECT 61.110 201.850 61.430 202.110 ;
        RECT 69.940 202.095 70.080 202.250 ;
        RECT 69.865 201.865 70.155 202.095 ;
        RECT 72.165 202.050 72.455 202.095 ;
        RECT 73.070 202.050 73.390 202.110 ;
        RECT 73.620 202.095 73.760 202.250 ;
        RECT 76.290 202.250 77.900 202.390 ;
        RECT 82.385 202.390 82.675 202.435 ;
        RECT 85.505 202.390 85.795 202.435 ;
        RECT 87.395 202.390 87.685 202.435 ;
        RECT 82.385 202.250 87.685 202.390 ;
        RECT 76.290 202.190 76.610 202.250 ;
        RECT 82.385 202.205 82.675 202.250 ;
        RECT 85.505 202.205 85.795 202.250 ;
        RECT 87.395 202.205 87.685 202.250 ;
        RECT 72.165 201.910 73.390 202.050 ;
        RECT 72.165 201.865 72.455 201.910 ;
        RECT 73.070 201.850 73.390 201.910 ;
        RECT 73.545 202.050 73.835 202.095 ;
        RECT 74.450 202.050 74.770 202.110 ;
        RECT 73.545 201.910 74.770 202.050 ;
        RECT 73.545 201.865 73.835 201.910 ;
        RECT 74.450 201.850 74.770 201.910 ;
        RECT 79.050 202.050 79.370 202.110 ;
        RECT 79.525 202.050 79.815 202.095 ;
        RECT 79.050 201.910 79.815 202.050 ;
        RECT 79.050 201.850 79.370 201.910 ;
        RECT 79.525 201.865 79.815 201.910 ;
        RECT 84.570 202.050 84.890 202.110 ;
        RECT 86.885 202.050 87.175 202.095 ;
        RECT 84.570 201.910 87.175 202.050 ;
        RECT 84.570 201.850 84.890 201.910 ;
        RECT 86.885 201.865 87.175 201.910 ;
        RECT 60.210 201.710 60.500 201.755 ;
        RECT 62.045 201.710 62.335 201.755 ;
        RECT 65.625 201.710 65.915 201.755 ;
        RECT 60.210 201.570 65.915 201.710 ;
        RECT 60.210 201.525 60.500 201.570 ;
        RECT 62.045 201.525 62.335 201.570 ;
        RECT 65.625 201.525 65.915 201.570 ;
        RECT 63.405 201.370 64.055 201.415 ;
        RECT 64.790 201.370 65.110 201.430 ;
        RECT 66.705 201.415 66.995 201.730 ;
        RECT 71.120 201.710 71.410 201.755 ;
        RECT 73.990 201.710 74.310 201.770 ;
        RECT 71.120 201.570 74.310 201.710 ;
        RECT 71.120 201.525 71.410 201.570 ;
        RECT 73.990 201.510 74.310 201.570 ;
        RECT 66.705 201.370 67.295 201.415 ;
        RECT 63.405 201.230 67.295 201.370 ;
        RECT 63.405 201.185 64.055 201.230 ;
        RECT 64.790 201.170 65.110 201.230 ;
        RECT 67.005 201.185 67.295 201.230 ;
        RECT 74.910 201.170 75.230 201.430 ;
        RECT 75.370 201.370 75.690 201.430 ;
        RECT 77.525 201.370 77.815 201.415 ;
        RECT 75.370 201.230 77.815 201.370 ;
        RECT 75.370 201.170 75.690 201.230 ;
        RECT 77.525 201.185 77.815 201.230 ;
        RECT 78.605 201.370 78.895 201.415 ;
        RECT 79.510 201.370 79.830 201.430 ;
        RECT 81.305 201.415 81.595 201.730 ;
        RECT 82.385 201.710 82.675 201.755 ;
        RECT 85.965 201.710 86.255 201.755 ;
        RECT 87.800 201.710 88.090 201.755 ;
        RECT 82.385 201.570 88.090 201.710 ;
        RECT 82.385 201.525 82.675 201.570 ;
        RECT 85.965 201.525 86.255 201.570 ;
        RECT 87.800 201.525 88.090 201.570 ;
        RECT 88.250 201.710 88.570 201.770 ;
        RECT 96.530 201.710 96.850 201.770 ;
        RECT 88.250 201.570 96.850 201.710 ;
        RECT 88.250 201.510 88.570 201.570 ;
        RECT 96.530 201.510 96.850 201.570 ;
        RECT 78.605 201.230 79.830 201.370 ;
        RECT 78.605 201.185 78.895 201.230 ;
        RECT 79.510 201.170 79.830 201.230 ;
        RECT 81.005 201.370 81.595 201.415 ;
        RECT 84.245 201.370 84.895 201.415 ;
        RECT 85.490 201.370 85.810 201.430 ;
        RECT 81.005 201.230 85.810 201.370 ;
        RECT 81.005 201.185 81.295 201.230 ;
        RECT 84.245 201.185 84.895 201.230 ;
        RECT 85.490 201.170 85.810 201.230 ;
        RECT 71.690 200.830 72.010 201.090 ;
        RECT 72.610 201.030 72.930 201.090 ;
        RECT 74.465 201.030 74.755 201.075 ;
        RECT 72.610 200.890 74.755 201.030 ;
        RECT 72.610 200.830 72.930 200.890 ;
        RECT 74.465 200.845 74.755 200.890 ;
        RECT 75.830 201.030 76.150 201.090 ;
        RECT 76.765 201.030 77.055 201.075 ;
        RECT 75.830 200.890 77.055 201.030 ;
        RECT 75.830 200.830 76.150 200.890 ;
        RECT 76.765 200.845 77.055 200.890 ;
        RECT 14.580 200.210 127.740 200.690 ;
        RECT 61.110 200.010 61.430 200.070 ;
        RECT 67.565 200.010 67.855 200.055 ;
        RECT 72.165 200.010 72.455 200.055 ;
        RECT 73.990 200.010 74.310 200.070 ;
        RECT 61.110 199.870 67.855 200.010 ;
        RECT 61.110 199.810 61.430 199.870 ;
        RECT 67.565 199.825 67.855 199.870 ;
        RECT 71.090 199.870 74.310 200.010 ;
        RECT 69.865 199.670 70.155 199.715 ;
        RECT 71.090 199.670 71.230 199.870 ;
        RECT 72.165 199.825 72.455 199.870 ;
        RECT 73.990 199.810 74.310 199.870 ;
        RECT 74.910 200.010 75.230 200.070 ;
        RECT 75.385 200.010 75.675 200.055 ;
        RECT 74.910 199.870 75.675 200.010 ;
        RECT 74.910 199.810 75.230 199.870 ;
        RECT 75.385 199.825 75.675 199.870 ;
        RECT 76.290 200.010 76.610 200.070 ;
        RECT 79.065 200.010 79.355 200.055 ;
        RECT 76.290 199.870 79.355 200.010 ;
        RECT 76.290 199.810 76.610 199.870 ;
        RECT 79.065 199.825 79.355 199.870 ;
        RECT 79.510 200.010 79.830 200.070 ;
        RECT 81.365 200.010 81.655 200.055 ;
        RECT 79.510 199.870 81.655 200.010 ;
        RECT 79.510 199.810 79.830 199.870 ;
        RECT 81.365 199.825 81.655 199.870 ;
        RECT 83.650 199.810 83.970 200.070 ;
        RECT 84.570 199.810 84.890 200.070 ;
        RECT 85.490 200.010 85.810 200.070 ;
        RECT 85.965 200.010 86.255 200.055 ;
        RECT 85.490 199.870 86.255 200.010 ;
        RECT 85.490 199.810 85.810 199.870 ;
        RECT 85.965 199.825 86.255 199.870 ;
        RECT 69.865 199.530 71.230 199.670 ;
        RECT 69.865 199.485 70.155 199.530 ;
        RECT 74.450 199.470 74.770 199.730 ;
        RECT 80.890 199.670 81.210 199.730 ;
        RECT 97.910 199.670 98.230 199.730 ;
        RECT 98.485 199.670 98.775 199.715 ;
        RECT 101.725 199.670 102.375 199.715 ;
        RECT 80.890 199.530 84.340 199.670 ;
        RECT 80.890 199.470 81.210 199.530 ;
        RECT 68.470 199.130 68.790 199.390 ;
        RECT 71.690 199.330 72.010 199.390 ;
        RECT 78.605 199.330 78.895 199.375 ;
        RECT 79.050 199.330 79.370 199.390 ;
        RECT 71.690 199.190 79.370 199.330 ;
        RECT 71.690 199.130 72.010 199.190 ;
        RECT 78.605 199.145 78.895 199.190 ;
        RECT 79.050 199.130 79.370 199.190 ;
        RECT 79.970 199.330 80.290 199.390 ;
        RECT 82.360 199.375 82.500 199.530 ;
        RECT 84.200 199.375 84.340 199.530 ;
        RECT 97.910 199.530 102.375 199.670 ;
        RECT 97.910 199.470 98.230 199.530 ;
        RECT 98.485 199.485 99.075 199.530 ;
        RECT 101.725 199.485 102.375 199.530 ;
        RECT 81.365 199.330 81.655 199.375 ;
        RECT 79.970 199.190 81.655 199.330 ;
        RECT 79.970 199.130 80.290 199.190 ;
        RECT 81.365 199.145 81.655 199.190 ;
        RECT 82.285 199.145 82.575 199.375 ;
        RECT 82.745 199.145 83.035 199.375 ;
        RECT 84.125 199.145 84.415 199.375 ;
        RECT 86.425 199.330 86.715 199.375 ;
        RECT 86.870 199.330 87.190 199.390 ;
        RECT 86.425 199.190 87.190 199.330 ;
        RECT 86.425 199.145 86.715 199.190 ;
        RECT 75.830 198.990 76.150 199.050 ;
        RECT 82.820 198.990 82.960 199.145 ;
        RECT 86.870 199.130 87.190 199.190 ;
        RECT 98.785 199.170 99.075 199.485 ;
        RECT 99.865 199.330 100.155 199.375 ;
        RECT 103.445 199.330 103.735 199.375 ;
        RECT 105.280 199.330 105.570 199.375 ;
        RECT 99.865 199.190 105.570 199.330 ;
        RECT 99.865 199.145 100.155 199.190 ;
        RECT 103.445 199.145 103.735 199.190 ;
        RECT 105.280 199.145 105.570 199.190 ;
        RECT 75.830 198.850 82.960 198.990 ;
        RECT 75.830 198.790 76.150 198.850 ;
        RECT 104.350 198.790 104.670 199.050 ;
        RECT 105.730 198.790 106.050 199.050 ;
        RECT 68.945 198.650 69.235 198.695 ;
        RECT 73.070 198.650 73.390 198.710 ;
        RECT 68.945 198.510 73.390 198.650 ;
        RECT 68.945 198.465 69.235 198.510 ;
        RECT 73.070 198.450 73.390 198.510 ;
        RECT 73.530 198.650 73.850 198.710 ;
        RECT 74.465 198.650 74.755 198.695 ;
        RECT 73.530 198.510 74.755 198.650 ;
        RECT 73.530 198.450 73.850 198.510 ;
        RECT 74.465 198.465 74.755 198.510 ;
        RECT 99.865 198.650 100.155 198.695 ;
        RECT 102.985 198.650 103.275 198.695 ;
        RECT 104.875 198.650 105.165 198.695 ;
        RECT 99.865 198.510 105.165 198.650 ;
        RECT 99.865 198.465 100.155 198.510 ;
        RECT 102.985 198.465 103.275 198.510 ;
        RECT 104.875 198.465 105.165 198.510 ;
        RECT 64.790 198.310 65.110 198.370 ;
        RECT 70.785 198.310 71.075 198.355 ;
        RECT 64.790 198.170 71.075 198.310 ;
        RECT 64.790 198.110 65.110 198.170 ;
        RECT 70.785 198.125 71.075 198.170 ;
        RECT 72.610 198.310 72.930 198.370 ;
        RECT 80.890 198.310 81.210 198.370 ;
        RECT 72.610 198.170 81.210 198.310 ;
        RECT 72.610 198.110 72.930 198.170 ;
        RECT 80.890 198.110 81.210 198.170 ;
        RECT 97.005 198.310 97.295 198.355 ;
        RECT 98.370 198.310 98.690 198.370 ;
        RECT 97.005 198.170 98.690 198.310 ;
        RECT 97.005 198.125 97.295 198.170 ;
        RECT 98.370 198.110 98.690 198.170 ;
        RECT 14.580 197.490 127.740 197.970 ;
        RECT 68.470 197.290 68.790 197.350 ;
        RECT 68.945 197.290 69.235 197.335 ;
        RECT 68.470 197.150 69.235 197.290 ;
        RECT 68.470 197.090 68.790 197.150 ;
        RECT 68.945 197.105 69.235 197.150 ;
        RECT 69.850 197.090 70.170 197.350 ;
        RECT 73.530 197.290 73.850 197.350 ;
        RECT 72.240 197.150 73.850 197.290 ;
        RECT 50.530 196.610 50.850 196.670 ;
        RECT 54.225 196.610 54.515 196.655 ;
        RECT 50.530 196.470 54.515 196.610 ;
        RECT 50.530 196.410 50.850 196.470 ;
        RECT 54.225 196.425 54.515 196.470 ;
        RECT 70.310 196.610 70.630 196.670 ;
        RECT 72.240 196.655 72.380 197.150 ;
        RECT 73.530 197.090 73.850 197.150 ;
        RECT 79.970 196.950 80.290 197.010 ;
        RECT 73.620 196.810 80.290 196.950 ;
        RECT 72.165 196.610 72.455 196.655 ;
        RECT 70.310 196.470 72.455 196.610 ;
        RECT 70.310 196.410 70.630 196.470 ;
        RECT 72.165 196.425 72.455 196.470 ;
        RECT 72.610 196.410 72.930 196.670 ;
        RECT 73.070 196.610 73.390 196.670 ;
        RECT 73.620 196.610 73.760 196.810 ;
        RECT 79.970 196.750 80.290 196.810 ;
        RECT 89.600 196.950 89.890 196.995 ;
        RECT 92.380 196.950 92.670 196.995 ;
        RECT 94.240 196.950 94.530 196.995 ;
        RECT 89.600 196.810 94.530 196.950 ;
        RECT 89.600 196.765 89.890 196.810 ;
        RECT 92.380 196.765 92.670 196.810 ;
        RECT 94.240 196.765 94.530 196.810 ;
        RECT 113.205 196.950 113.495 196.995 ;
        RECT 116.325 196.950 116.615 196.995 ;
        RECT 118.215 196.950 118.505 196.995 ;
        RECT 113.205 196.810 118.505 196.950 ;
        RECT 113.205 196.765 113.495 196.810 ;
        RECT 116.325 196.765 116.615 196.810 ;
        RECT 118.215 196.765 118.505 196.810 ;
        RECT 73.070 196.470 73.760 196.610 ;
        RECT 92.865 196.610 93.155 196.655 ;
        RECT 93.770 196.610 94.090 196.670 ;
        RECT 92.865 196.470 94.090 196.610 ;
        RECT 73.070 196.410 73.390 196.470 ;
        RECT 92.865 196.425 93.155 196.470 ;
        RECT 93.770 196.410 94.090 196.470 ;
        RECT 49.150 196.270 49.470 196.330 ;
        RECT 53.765 196.270 54.055 196.315 ;
        RECT 49.150 196.130 54.055 196.270 ;
        RECT 49.150 196.070 49.470 196.130 ;
        RECT 53.765 196.085 54.055 196.130 ;
        RECT 68.930 196.270 69.250 196.330 ;
        RECT 73.545 196.270 73.835 196.315 ;
        RECT 74.450 196.270 74.770 196.330 ;
        RECT 68.930 196.130 74.770 196.270 ;
        RECT 68.930 196.070 69.250 196.130 ;
        RECT 73.545 196.085 73.835 196.130 ;
        RECT 74.450 196.070 74.770 196.130 ;
        RECT 89.600 196.270 89.890 196.315 ;
        RECT 94.705 196.270 94.995 196.315 ;
        RECT 96.530 196.270 96.850 196.330 ;
        RECT 89.600 196.130 92.135 196.270 ;
        RECT 89.600 196.085 89.890 196.130 ;
        RECT 70.785 195.930 71.075 195.975 ;
        RECT 71.690 195.930 72.010 195.990 ;
        RECT 75.370 195.930 75.690 195.990 ;
        RECT 70.785 195.790 75.690 195.930 ;
        RECT 70.785 195.745 71.075 195.790 ;
        RECT 71.690 195.730 72.010 195.790 ;
        RECT 75.370 195.730 75.690 195.790 ;
        RECT 87.740 195.930 88.030 195.975 ;
        RECT 90.090 195.930 90.410 195.990 ;
        RECT 91.920 195.975 92.135 196.130 ;
        RECT 94.705 196.130 96.850 196.270 ;
        RECT 94.705 196.085 94.995 196.130 ;
        RECT 96.530 196.070 96.850 196.130 ;
        RECT 98.370 196.070 98.690 196.330 ;
        RECT 112.125 195.975 112.415 196.290 ;
        RECT 113.205 196.270 113.495 196.315 ;
        RECT 116.785 196.270 117.075 196.315 ;
        RECT 118.620 196.270 118.910 196.315 ;
        RECT 113.205 196.130 118.910 196.270 ;
        RECT 113.205 196.085 113.495 196.130 ;
        RECT 116.785 196.085 117.075 196.130 ;
        RECT 118.620 196.085 118.910 196.130 ;
        RECT 119.085 196.085 119.375 196.315 ;
        RECT 115.390 195.975 115.710 195.990 ;
        RECT 91.000 195.930 91.290 195.975 ;
        RECT 87.740 195.790 91.290 195.930 ;
        RECT 87.740 195.745 88.030 195.790 ;
        RECT 90.090 195.730 90.410 195.790 ;
        RECT 91.000 195.745 91.290 195.790 ;
        RECT 91.920 195.930 92.210 195.975 ;
        RECT 93.780 195.930 94.070 195.975 ;
        RECT 91.920 195.790 94.070 195.930 ;
        RECT 91.920 195.745 92.210 195.790 ;
        RECT 93.780 195.745 94.070 195.790 ;
        RECT 111.825 195.930 112.415 195.975 ;
        RECT 115.065 195.930 115.715 195.975 ;
        RECT 111.825 195.790 115.715 195.930 ;
        RECT 111.825 195.745 112.115 195.790 ;
        RECT 115.065 195.745 115.715 195.790 ;
        RECT 115.390 195.730 115.710 195.745 ;
        RECT 117.690 195.730 118.010 195.990 ;
        RECT 118.150 195.930 118.470 195.990 ;
        RECT 119.160 195.930 119.300 196.085 ;
        RECT 118.150 195.790 119.300 195.930 ;
        RECT 118.150 195.730 118.470 195.790 ;
        RECT 53.290 195.390 53.610 195.650 ;
        RECT 57.445 195.590 57.735 195.635 ;
        RECT 57.890 195.590 58.210 195.650 ;
        RECT 85.490 195.635 85.810 195.650 ;
        RECT 57.445 195.450 58.210 195.590 ;
        RECT 57.445 195.405 57.735 195.450 ;
        RECT 57.890 195.390 58.210 195.450 ;
        RECT 69.785 195.590 70.075 195.635 ;
        RECT 71.245 195.590 71.535 195.635 ;
        RECT 69.785 195.450 71.535 195.590 ;
        RECT 69.785 195.405 70.075 195.450 ;
        RECT 71.245 195.405 71.535 195.450 ;
        RECT 85.490 195.405 86.025 195.635 ;
        RECT 85.490 195.390 85.810 195.405 ;
        RECT 101.130 195.390 101.450 195.650 ;
        RECT 108.950 195.590 109.270 195.650 ;
        RECT 110.345 195.590 110.635 195.635 ;
        RECT 108.950 195.450 110.635 195.590 ;
        RECT 108.950 195.390 109.270 195.450 ;
        RECT 110.345 195.405 110.635 195.450 ;
        RECT 14.580 194.770 127.740 195.250 ;
        RECT 50.530 194.570 50.850 194.630 ;
        RECT 57.905 194.570 58.195 194.615 ;
        RECT 50.530 194.430 58.195 194.570 ;
        RECT 50.530 194.370 50.850 194.430 ;
        RECT 57.905 194.385 58.195 194.430 ;
        RECT 71.690 194.370 72.010 194.630 ;
        RECT 85.490 194.570 85.810 194.630 ;
        RECT 85.965 194.570 86.255 194.615 ;
        RECT 72.240 194.430 85.260 194.570 ;
        RECT 49.150 194.230 49.470 194.290 ;
        RECT 53.290 194.275 53.610 194.290 ;
        RECT 48.780 194.090 49.470 194.230 ;
        RECT 45.930 193.890 46.250 193.950 ;
        RECT 48.780 193.935 48.920 194.090 ;
        RECT 49.150 194.030 49.470 194.090 ;
        RECT 52.825 194.230 53.610 194.275 ;
        RECT 56.425 194.230 56.715 194.275 ;
        RECT 72.240 194.230 72.380 194.430 ;
        RECT 52.825 194.090 56.715 194.230 ;
        RECT 52.825 194.045 53.610 194.090 ;
        RECT 53.290 194.030 53.610 194.045 ;
        RECT 56.125 194.045 56.715 194.090 ;
        RECT 66.260 194.090 72.380 194.230 ;
        RECT 72.610 194.230 72.930 194.290 ;
        RECT 85.120 194.230 85.260 194.430 ;
        RECT 85.490 194.430 86.255 194.570 ;
        RECT 85.490 194.370 85.810 194.430 ;
        RECT 85.965 194.385 86.255 194.430 ;
        RECT 89.645 194.570 89.935 194.615 ;
        RECT 90.090 194.570 90.410 194.630 ;
        RECT 89.645 194.430 90.410 194.570 ;
        RECT 89.645 194.385 89.935 194.430 ;
        RECT 90.090 194.370 90.410 194.430 ;
        RECT 93.785 194.570 94.075 194.615 ;
        RECT 97.910 194.570 98.230 194.630 ;
        RECT 93.785 194.430 98.230 194.570 ;
        RECT 93.785 194.385 94.075 194.430 ;
        RECT 97.910 194.370 98.230 194.430 ;
        RECT 112.185 194.570 112.475 194.615 ;
        RECT 112.630 194.570 112.950 194.630 ;
        RECT 112.185 194.430 112.950 194.570 ;
        RECT 112.185 194.385 112.475 194.430 ;
        RECT 112.630 194.370 112.950 194.430 ;
        RECT 115.390 194.370 115.710 194.630 ;
        RECT 86.870 194.230 87.190 194.290 ;
        RECT 96.530 194.230 96.850 194.290 ;
        RECT 103.445 194.230 103.735 194.275 ;
        RECT 105.730 194.230 106.050 194.290 ;
        RECT 118.150 194.230 118.470 194.290 ;
        RECT 72.610 194.090 75.140 194.230 ;
        RECT 85.120 194.090 95.380 194.230 ;
        RECT 48.705 193.890 48.995 193.935 ;
        RECT 45.930 193.750 48.995 193.890 ;
        RECT 45.930 193.690 46.250 193.750 ;
        RECT 48.705 193.705 48.995 193.750 ;
        RECT 49.630 193.890 49.920 193.935 ;
        RECT 51.465 193.890 51.755 193.935 ;
        RECT 55.045 193.890 55.335 193.935 ;
        RECT 49.630 193.750 55.335 193.890 ;
        RECT 49.630 193.705 49.920 193.750 ;
        RECT 51.465 193.705 51.755 193.750 ;
        RECT 55.045 193.705 55.335 193.750 ;
        RECT 56.125 193.730 56.415 194.045 ;
        RECT 66.260 193.950 66.400 194.090 ;
        RECT 72.610 194.030 72.930 194.090 ;
        RECT 66.170 193.690 66.490 193.950 ;
        RECT 68.930 193.690 69.250 193.950 ;
        RECT 73.070 193.690 73.390 193.950 ;
        RECT 75.000 193.935 75.140 194.090 ;
        RECT 86.870 194.030 87.190 194.090 ;
        RECT 74.925 193.890 75.215 193.935 ;
        RECT 76.290 193.890 76.610 193.950 ;
        RECT 74.925 193.750 76.610 193.890 ;
        RECT 74.925 193.705 75.215 193.750 ;
        RECT 76.290 193.690 76.610 193.750 ;
        RECT 85.950 193.890 86.270 193.950 ;
        RECT 86.425 193.890 86.715 193.935 ;
        RECT 85.950 193.750 86.715 193.890 ;
        RECT 85.950 193.690 86.270 193.750 ;
        RECT 86.425 193.705 86.715 193.750 ;
        RECT 90.090 193.690 90.410 193.950 ;
        RECT 93.400 193.935 93.540 194.090 ;
        RECT 93.325 193.705 93.615 193.935 ;
        RECT 94.690 193.690 95.010 193.950 ;
        RECT 95.240 193.890 95.380 194.090 ;
        RECT 96.530 194.090 118.470 194.230 ;
        RECT 96.530 194.030 96.850 194.090 ;
        RECT 103.445 194.045 103.735 194.090 ;
        RECT 105.730 194.030 106.050 194.090 ;
        RECT 118.150 194.030 118.470 194.090 ;
        RECT 108.965 193.890 109.255 193.935 ;
        RECT 115.850 193.890 116.170 193.950 ;
        RECT 95.240 193.750 116.170 193.890 ;
        RECT 108.965 193.705 109.255 193.750 ;
        RECT 115.850 193.690 116.170 193.750 ;
        RECT 49.150 193.350 49.470 193.610 ;
        RECT 50.530 193.350 50.850 193.610 ;
        RECT 70.325 193.550 70.615 193.595 ;
        RECT 70.325 193.410 72.380 193.550 ;
        RECT 70.325 193.365 70.615 193.410 ;
        RECT 72.240 193.255 72.380 193.410 ;
        RECT 85.030 193.350 85.350 193.610 ;
        RECT 108.030 193.550 108.350 193.610 ;
        RECT 110.790 193.550 111.110 193.610 ;
        RECT 108.030 193.410 111.110 193.550 ;
        RECT 108.030 193.350 108.350 193.410 ;
        RECT 110.790 193.350 111.110 193.410 ;
        RECT 111.725 193.365 112.015 193.595 ;
        RECT 50.035 193.210 50.325 193.255 ;
        RECT 51.925 193.210 52.215 193.255 ;
        RECT 55.045 193.210 55.335 193.255 ;
        RECT 50.035 193.070 55.335 193.210 ;
        RECT 50.035 193.025 50.325 193.070 ;
        RECT 51.925 193.025 52.215 193.070 ;
        RECT 55.045 193.025 55.335 193.070 ;
        RECT 72.165 193.025 72.455 193.255 ;
        RECT 111.800 193.210 111.940 193.365 ;
        RECT 112.170 193.210 112.490 193.270 ;
        RECT 111.800 193.070 112.490 193.210 ;
        RECT 112.170 193.010 112.490 193.070 ;
        RECT 48.245 192.870 48.535 192.915 ;
        RECT 54.210 192.870 54.530 192.930 ;
        RECT 48.245 192.730 54.530 192.870 ;
        RECT 48.245 192.685 48.535 192.730 ;
        RECT 54.210 192.670 54.530 192.730 ;
        RECT 65.710 192.670 66.030 192.930 ;
        RECT 70.310 192.670 70.630 192.930 ;
        RECT 72.610 192.870 72.930 192.930 ;
        RECT 73.085 192.870 73.375 192.915 ;
        RECT 72.610 192.730 73.375 192.870 ;
        RECT 72.610 192.670 72.930 192.730 ;
        RECT 73.085 192.685 73.375 192.730 ;
        RECT 88.265 192.870 88.555 192.915 ;
        RECT 91.010 192.870 91.330 192.930 ;
        RECT 88.265 192.730 91.330 192.870 ;
        RECT 88.265 192.685 88.555 192.730 ;
        RECT 91.010 192.670 91.330 192.730 ;
        RECT 109.410 192.670 109.730 192.930 ;
        RECT 114.025 192.870 114.315 192.915 ;
        RECT 119.070 192.870 119.390 192.930 ;
        RECT 114.025 192.730 119.390 192.870 ;
        RECT 114.025 192.685 114.315 192.730 ;
        RECT 119.070 192.670 119.390 192.730 ;
        RECT 14.580 192.050 127.740 192.530 ;
        RECT 50.530 191.850 50.850 191.910 ;
        RECT 51.005 191.850 51.295 191.895 ;
        RECT 50.530 191.710 51.295 191.850 ;
        RECT 50.530 191.650 50.850 191.710 ;
        RECT 51.005 191.665 51.295 191.710 ;
        RECT 85.490 191.850 85.810 191.910 ;
        RECT 85.490 191.710 93.540 191.850 ;
        RECT 85.490 191.650 85.810 191.710 ;
        RECT 40.380 191.510 40.670 191.555 ;
        RECT 43.160 191.510 43.450 191.555 ;
        RECT 45.020 191.510 45.310 191.555 ;
        RECT 40.380 191.370 45.310 191.510 ;
        RECT 40.380 191.325 40.670 191.370 ;
        RECT 43.160 191.325 43.450 191.370 ;
        RECT 45.020 191.325 45.310 191.370 ;
        RECT 49.625 191.325 49.915 191.555 ;
        RECT 55.245 191.510 55.535 191.555 ;
        RECT 58.365 191.510 58.655 191.555 ;
        RECT 60.255 191.510 60.545 191.555 ;
        RECT 55.245 191.370 60.545 191.510 ;
        RECT 55.245 191.325 55.535 191.370 ;
        RECT 58.365 191.325 58.655 191.370 ;
        RECT 60.255 191.325 60.545 191.370 ;
        RECT 36.515 191.170 36.805 191.215 ;
        RECT 41.330 191.170 41.650 191.230 ;
        RECT 36.515 191.030 46.160 191.170 ;
        RECT 36.515 190.985 36.805 191.030 ;
        RECT 41.330 190.970 41.650 191.030 ;
        RECT 40.380 190.830 40.670 190.875 ;
        RECT 43.645 190.830 43.935 190.875 ;
        RECT 45.010 190.830 45.330 190.890 ;
        RECT 40.380 190.690 42.915 190.830 ;
        RECT 40.380 190.645 40.670 190.690 ;
        RECT 38.520 190.490 38.810 190.535 ;
        RECT 39.030 190.490 39.350 190.550 ;
        RECT 42.700 190.535 42.915 190.690 ;
        RECT 43.645 190.690 45.330 190.830 ;
        RECT 43.645 190.645 43.935 190.690 ;
        RECT 45.010 190.630 45.330 190.690 ;
        RECT 45.485 190.645 45.775 190.875 ;
        RECT 46.020 190.830 46.160 191.030 ;
        RECT 46.390 190.970 46.710 191.230 ;
        RECT 47.785 190.830 48.075 190.875 ;
        RECT 46.020 190.690 48.075 190.830 ;
        RECT 49.700 190.830 49.840 191.325 ;
        RECT 63.870 191.310 64.190 191.570 ;
        RECT 64.905 191.510 65.195 191.555 ;
        RECT 68.025 191.510 68.315 191.555 ;
        RECT 69.915 191.510 70.205 191.555 ;
        RECT 76.765 191.510 77.055 191.555 ;
        RECT 64.905 191.370 70.205 191.510 ;
        RECT 64.905 191.325 65.195 191.370 ;
        RECT 68.025 191.325 68.315 191.370 ;
        RECT 69.915 191.325 70.205 191.370 ;
        RECT 73.620 191.370 77.055 191.510 ;
        RECT 52.370 190.970 52.690 191.230 ;
        RECT 59.270 191.170 59.590 191.230 ;
        RECT 61.125 191.170 61.415 191.215 ;
        RECT 63.960 191.170 64.100 191.310 ;
        RECT 70.785 191.170 71.075 191.215 ;
        RECT 59.270 191.030 71.075 191.170 ;
        RECT 59.270 190.970 59.590 191.030 ;
        RECT 61.125 190.985 61.415 191.030 ;
        RECT 70.785 190.985 71.075 191.030 ;
        RECT 71.230 191.170 71.550 191.230 ;
        RECT 73.620 191.215 73.760 191.370 ;
        RECT 76.765 191.325 77.055 191.370 ;
        RECT 87.300 191.510 87.590 191.555 ;
        RECT 90.080 191.510 90.370 191.555 ;
        RECT 91.940 191.510 92.230 191.555 ;
        RECT 87.300 191.370 92.230 191.510 ;
        RECT 93.400 191.510 93.540 191.710 ;
        RECT 93.770 191.650 94.090 191.910 ;
        RECT 102.985 191.850 103.275 191.895 ;
        RECT 104.350 191.850 104.670 191.910 ;
        RECT 112.630 191.850 112.950 191.910 ;
        RECT 102.985 191.710 104.670 191.850 ;
        RECT 102.985 191.665 103.275 191.710 ;
        RECT 104.350 191.650 104.670 191.710 ;
        RECT 108.580 191.710 112.950 191.850 ;
        RECT 108.030 191.510 108.350 191.570 ;
        RECT 93.400 191.370 97.220 191.510 ;
        RECT 87.300 191.325 87.590 191.370 ;
        RECT 90.080 191.325 90.370 191.370 ;
        RECT 91.940 191.325 92.230 191.370 ;
        RECT 73.545 191.170 73.835 191.215 ;
        RECT 71.230 191.030 73.835 191.170 ;
        RECT 71.230 190.970 71.550 191.030 ;
        RECT 73.545 190.985 73.835 191.030 ;
        RECT 78.145 191.170 78.435 191.215 ;
        RECT 79.970 191.170 80.290 191.230 ;
        RECT 78.145 191.030 80.290 191.170 ;
        RECT 78.145 190.985 78.435 191.030 ;
        RECT 79.970 190.970 80.290 191.030 ;
        RECT 92.405 191.170 92.695 191.215 ;
        RECT 93.770 191.170 94.090 191.230 ;
        RECT 92.405 191.030 96.760 191.170 ;
        RECT 92.405 190.985 92.695 191.030 ;
        RECT 93.770 190.970 94.090 191.030 ;
        RECT 96.620 190.890 96.760 191.030 ;
        RECT 51.925 190.830 52.215 190.875 ;
        RECT 54.210 190.850 54.530 190.890 ;
        RECT 49.700 190.690 52.215 190.830 ;
        RECT 47.785 190.645 48.075 190.690 ;
        RECT 51.925 190.645 52.215 190.690 ;
        RECT 41.780 190.490 42.070 190.535 ;
        RECT 38.520 190.350 42.070 190.490 ;
        RECT 38.520 190.305 38.810 190.350 ;
        RECT 39.030 190.290 39.350 190.350 ;
        RECT 41.780 190.305 42.070 190.350 ;
        RECT 42.700 190.490 42.990 190.535 ;
        RECT 44.560 190.490 44.850 190.535 ;
        RECT 42.700 190.350 44.850 190.490 ;
        RECT 45.560 190.490 45.700 190.645 ;
        RECT 54.165 190.630 54.530 190.850 ;
        RECT 55.245 190.830 55.535 190.875 ;
        RECT 58.825 190.830 59.115 190.875 ;
        RECT 60.660 190.830 60.950 190.875 ;
        RECT 55.245 190.690 60.950 190.830 ;
        RECT 55.245 190.645 55.535 190.690 ;
        RECT 58.825 190.645 59.115 190.690 ;
        RECT 60.660 190.645 60.950 190.690 ;
        RECT 49.150 190.490 49.470 190.550 ;
        RECT 54.165 190.535 54.455 190.630 ;
        RECT 45.560 190.350 49.470 190.490 ;
        RECT 42.700 190.305 42.990 190.350 ;
        RECT 44.560 190.305 44.850 190.350 ;
        RECT 49.150 190.290 49.470 190.350 ;
        RECT 53.865 190.490 54.455 190.535 ;
        RECT 57.105 190.490 57.755 190.535 ;
        RECT 53.865 190.350 57.755 190.490 ;
        RECT 53.865 190.305 54.155 190.350 ;
        RECT 57.105 190.305 57.755 190.350 ;
        RECT 59.745 190.490 60.035 190.535 ;
        RECT 60.190 190.490 60.510 190.550 ;
        RECT 63.825 190.535 64.115 190.850 ;
        RECT 64.905 190.830 65.195 190.875 ;
        RECT 68.485 190.830 68.775 190.875 ;
        RECT 70.320 190.830 70.610 190.875 ;
        RECT 64.905 190.690 70.610 190.830 ;
        RECT 64.905 190.645 65.195 190.690 ;
        RECT 68.485 190.645 68.775 190.690 ;
        RECT 70.320 190.645 70.610 190.690 ;
        RECT 73.070 190.630 73.390 190.890 ;
        RECT 74.450 190.830 74.770 190.890 ;
        RECT 76.305 190.830 76.595 190.875 ;
        RECT 74.450 190.690 76.595 190.830 ;
        RECT 74.450 190.630 74.770 190.690 ;
        RECT 76.305 190.645 76.595 190.690 ;
        RECT 87.300 190.830 87.590 190.875 ;
        RECT 87.300 190.690 89.835 190.830 ;
        RECT 87.300 190.645 87.590 190.690 ;
        RECT 59.745 190.350 60.510 190.490 ;
        RECT 59.745 190.305 60.035 190.350 ;
        RECT 60.190 190.290 60.510 190.350 ;
        RECT 63.525 190.490 64.115 190.535 ;
        RECT 65.710 190.490 66.030 190.550 ;
        RECT 66.765 190.490 67.415 190.535 ;
        RECT 63.525 190.350 67.415 190.490 ;
        RECT 63.525 190.305 63.815 190.350 ;
        RECT 65.710 190.290 66.030 190.350 ;
        RECT 66.765 190.305 67.415 190.350 ;
        RECT 69.405 190.490 69.695 190.535 ;
        RECT 73.530 190.490 73.850 190.550 ;
        RECT 76.765 190.490 77.055 190.535 ;
        RECT 69.405 190.350 71.460 190.490 ;
        RECT 69.405 190.305 69.695 190.350 ;
        RECT 47.325 190.150 47.615 190.195 ;
        RECT 57.890 190.150 58.210 190.210 ;
        RECT 47.325 190.010 58.210 190.150 ;
        RECT 47.325 189.965 47.615 190.010 ;
        RECT 57.890 189.950 58.210 190.010 ;
        RECT 62.030 189.950 62.350 190.210 ;
        RECT 66.170 190.150 66.490 190.210 ;
        RECT 69.850 190.150 70.170 190.210 ;
        RECT 71.320 190.195 71.460 190.350 ;
        RECT 73.530 190.350 77.055 190.490 ;
        RECT 73.530 190.290 73.850 190.350 ;
        RECT 76.765 190.305 77.055 190.350 ;
        RECT 85.440 190.490 85.730 190.535 ;
        RECT 87.790 190.490 88.110 190.550 ;
        RECT 89.620 190.535 89.835 190.690 ;
        RECT 90.550 190.630 90.870 190.890 ;
        RECT 91.010 190.830 91.330 190.890 ;
        RECT 92.865 190.830 93.155 190.875 ;
        RECT 91.010 190.690 93.155 190.830 ;
        RECT 91.010 190.630 91.330 190.690 ;
        RECT 92.865 190.645 93.155 190.690 ;
        RECT 96.530 190.630 96.850 190.890 ;
        RECT 97.080 190.830 97.220 191.370 ;
        RECT 98.000 191.370 108.350 191.510 ;
        RECT 98.000 191.230 98.140 191.370 ;
        RECT 97.910 190.970 98.230 191.230 ;
        RECT 98.845 191.170 99.135 191.215 ;
        RECT 101.130 191.170 101.450 191.230 ;
        RECT 105.360 191.215 105.500 191.370 ;
        RECT 108.030 191.310 108.350 191.370 ;
        RECT 98.845 191.030 102.740 191.170 ;
        RECT 98.845 190.985 99.135 191.030 ;
        RECT 101.130 190.970 101.450 191.030 ;
        RECT 99.305 190.830 99.595 190.875 ;
        RECT 102.065 190.830 102.355 190.875 ;
        RECT 97.080 190.690 99.595 190.830 ;
        RECT 99.305 190.645 99.595 190.690 ;
        RECT 101.220 190.690 102.355 190.830 ;
        RECT 102.600 190.830 102.740 191.030 ;
        RECT 105.285 190.985 105.575 191.215 ;
        RECT 106.190 191.170 106.510 191.230 ;
        RECT 108.580 191.170 108.720 191.710 ;
        RECT 112.630 191.650 112.950 191.710 ;
        RECT 117.690 191.850 118.010 191.910 ;
        RECT 118.165 191.850 118.455 191.895 ;
        RECT 117.690 191.710 118.455 191.850 ;
        RECT 117.690 191.650 118.010 191.710 ;
        RECT 118.165 191.665 118.455 191.710 ;
        RECT 111.825 191.510 112.115 191.555 ;
        RECT 114.945 191.510 115.235 191.555 ;
        RECT 116.835 191.510 117.125 191.555 ;
        RECT 111.825 191.370 117.125 191.510 ;
        RECT 111.825 191.325 112.115 191.370 ;
        RECT 114.945 191.325 115.235 191.370 ;
        RECT 116.835 191.325 117.125 191.370 ;
        RECT 106.190 191.030 108.720 191.170 ;
        RECT 108.965 191.170 109.255 191.215 ;
        RECT 109.870 191.170 110.190 191.230 ;
        RECT 108.965 191.030 110.190 191.170 ;
        RECT 106.190 190.970 106.510 191.030 ;
        RECT 108.965 190.985 109.255 191.030 ;
        RECT 109.870 190.970 110.190 191.030 ;
        RECT 106.665 190.830 106.955 190.875 ;
        RECT 102.600 190.690 106.955 190.830 ;
        RECT 88.700 190.490 88.990 190.535 ;
        RECT 85.440 190.350 88.990 190.490 ;
        RECT 85.440 190.305 85.730 190.350 ;
        RECT 87.790 190.290 88.110 190.350 ;
        RECT 88.700 190.305 88.990 190.350 ;
        RECT 89.620 190.490 89.910 190.535 ;
        RECT 91.480 190.490 91.770 190.535 ;
        RECT 89.620 190.350 91.770 190.490 ;
        RECT 89.620 190.305 89.910 190.350 ;
        RECT 91.480 190.305 91.770 190.350 ;
        RECT 66.170 190.010 70.170 190.150 ;
        RECT 66.170 189.950 66.490 190.010 ;
        RECT 69.850 189.950 70.170 190.010 ;
        RECT 71.245 189.965 71.535 190.195 ;
        RECT 76.290 190.150 76.610 190.210 ;
        RECT 77.225 190.150 77.515 190.195 ;
        RECT 76.290 190.010 77.515 190.150 ;
        RECT 76.290 189.950 76.610 190.010 ;
        RECT 77.225 189.965 77.515 190.010 ;
        RECT 83.435 190.150 83.725 190.195 ;
        RECT 85.950 190.150 86.270 190.210 ;
        RECT 101.220 190.195 101.360 190.690 ;
        RECT 102.065 190.645 102.355 190.690 ;
        RECT 106.665 190.645 106.955 190.690 ;
        RECT 109.410 190.490 109.730 190.550 ;
        RECT 110.745 190.535 111.035 190.850 ;
        RECT 111.825 190.830 112.115 190.875 ;
        RECT 115.405 190.830 115.695 190.875 ;
        RECT 117.240 190.830 117.530 190.875 ;
        RECT 111.825 190.690 117.530 190.830 ;
        RECT 111.825 190.645 112.115 190.690 ;
        RECT 115.405 190.645 115.695 190.690 ;
        RECT 117.240 190.645 117.530 190.690 ;
        RECT 117.705 190.830 117.995 190.875 ;
        RECT 118.150 190.830 118.470 190.890 ;
        RECT 117.705 190.690 118.470 190.830 ;
        RECT 117.705 190.645 117.995 190.690 ;
        RECT 118.150 190.630 118.470 190.690 ;
        RECT 119.070 190.630 119.390 190.890 ;
        RECT 110.445 190.490 111.035 190.535 ;
        RECT 113.685 190.490 114.335 190.535 ;
        RECT 109.410 190.350 114.335 190.490 ;
        RECT 109.410 190.290 109.730 190.350 ;
        RECT 110.445 190.305 110.735 190.350 ;
        RECT 113.685 190.305 114.335 190.350 ;
        RECT 116.310 190.290 116.630 190.550 ;
        RECT 83.435 190.010 86.270 190.150 ;
        RECT 83.435 189.965 83.725 190.010 ;
        RECT 85.950 189.950 86.270 190.010 ;
        RECT 101.145 189.965 101.435 190.195 ;
        RECT 108.505 190.150 108.795 190.195 ;
        RECT 113.090 190.150 113.410 190.210 ;
        RECT 108.505 190.010 113.410 190.150 ;
        RECT 108.505 189.965 108.795 190.010 ;
        RECT 113.090 189.950 113.410 190.010 ;
        RECT 14.580 189.330 127.740 189.810 ;
        RECT 57.890 188.930 58.210 189.190 ;
        RECT 59.745 188.945 60.035 189.175 ;
        RECT 36.285 188.790 36.575 188.835 ;
        RECT 39.145 188.790 39.435 188.835 ;
        RECT 42.385 188.790 43.035 188.835 ;
        RECT 36.285 188.650 43.035 188.790 ;
        RECT 36.285 188.605 36.575 188.650 ;
        RECT 39.145 188.605 39.735 188.650 ;
        RECT 42.385 188.605 43.035 188.650 ;
        RECT 30.305 188.450 30.595 188.495 ;
        RECT 35.825 188.450 36.115 188.495 ;
        RECT 30.305 188.310 36.500 188.450 ;
        RECT 30.305 188.265 30.595 188.310 ;
        RECT 35.825 188.265 36.115 188.310 ;
        RECT 36.360 188.170 36.500 188.310 ;
        RECT 39.445 188.290 39.735 188.605 ;
        RECT 40.525 188.450 40.815 188.495 ;
        RECT 44.105 188.450 44.395 188.495 ;
        RECT 45.940 188.450 46.230 188.495 ;
        RECT 40.525 188.310 46.230 188.450 ;
        RECT 40.525 188.265 40.815 188.310 ;
        RECT 44.105 188.265 44.395 188.310 ;
        RECT 45.940 188.265 46.230 188.310 ;
        RECT 55.590 188.250 55.910 188.510 ;
        RECT 56.510 188.450 56.830 188.510 ;
        RECT 57.445 188.450 57.735 188.495 ;
        RECT 56.510 188.310 57.735 188.450 ;
        RECT 59.820 188.450 59.960 188.945 ;
        RECT 60.190 188.930 60.510 189.190 ;
        RECT 67.105 189.130 67.395 189.175 ;
        RECT 73.070 189.130 73.390 189.190 ;
        RECT 67.105 188.990 73.390 189.130 ;
        RECT 67.105 188.945 67.395 188.990 ;
        RECT 73.070 188.930 73.390 188.990 ;
        RECT 87.345 189.130 87.635 189.175 ;
        RECT 87.790 189.130 88.110 189.190 ;
        RECT 87.345 188.990 88.110 189.130 ;
        RECT 87.345 188.945 87.635 188.990 ;
        RECT 87.790 188.930 88.110 188.990 ;
        RECT 90.105 189.130 90.395 189.175 ;
        RECT 90.550 189.130 90.870 189.190 ;
        RECT 90.105 188.990 90.870 189.130 ;
        RECT 90.105 188.945 90.395 188.990 ;
        RECT 90.550 188.930 90.870 188.990 ;
        RECT 106.190 189.130 106.510 189.190 ;
        RECT 107.125 189.130 107.415 189.175 ;
        RECT 106.190 188.990 107.415 189.130 ;
        RECT 106.190 188.930 106.510 188.990 ;
        RECT 107.125 188.945 107.415 188.990 ;
        RECT 114.025 189.130 114.315 189.175 ;
        RECT 116.310 189.130 116.630 189.190 ;
        RECT 114.025 188.990 116.630 189.130 ;
        RECT 114.025 188.945 114.315 188.990 ;
        RECT 116.310 188.930 116.630 188.990 ;
        RECT 99.405 188.790 99.695 188.835 ;
        RECT 100.210 188.790 100.530 188.850 ;
        RECT 102.645 188.790 103.295 188.835 ;
        RECT 99.405 188.650 103.295 188.790 ;
        RECT 99.405 188.605 99.995 188.650 ;
        RECT 61.125 188.450 61.415 188.495 ;
        RECT 59.820 188.310 61.415 188.450 ;
        RECT 56.510 188.250 56.830 188.310 ;
        RECT 57.445 188.265 57.735 188.310 ;
        RECT 61.125 188.265 61.415 188.310 ;
        RECT 87.805 188.265 88.095 188.495 ;
        RECT 28.450 188.110 28.770 188.170 ;
        RECT 29.845 188.110 30.135 188.155 ;
        RECT 28.450 187.970 30.135 188.110 ;
        RECT 28.450 187.910 28.770 187.970 ;
        RECT 29.845 187.925 30.135 187.970 ;
        RECT 36.270 187.910 36.590 188.170 ;
        RECT 44.550 188.110 44.870 188.170 ;
        RECT 46.405 188.110 46.695 188.155 ;
        RECT 44.550 187.970 46.695 188.110 ;
        RECT 44.550 187.910 44.870 187.970 ;
        RECT 46.405 187.925 46.695 187.970 ;
        RECT 46.850 188.110 47.170 188.170 ;
        RECT 56.985 188.110 57.275 188.155 ;
        RECT 46.850 187.970 57.275 188.110 ;
        RECT 40.525 187.770 40.815 187.815 ;
        RECT 43.645 187.770 43.935 187.815 ;
        RECT 45.535 187.770 45.825 187.815 ;
        RECT 40.525 187.630 45.825 187.770 ;
        RECT 46.480 187.770 46.620 187.925 ;
        RECT 46.850 187.910 47.170 187.970 ;
        RECT 56.985 187.925 57.275 187.970 ;
        RECT 62.030 188.110 62.350 188.170 ;
        RECT 64.345 188.110 64.635 188.155 ;
        RECT 65.710 188.110 66.030 188.170 ;
        RECT 72.150 188.110 72.470 188.170 ;
        RECT 62.030 187.970 72.470 188.110 ;
        RECT 87.880 188.110 88.020 188.265 ;
        RECT 89.170 188.250 89.490 188.510 ;
        RECT 99.705 188.290 99.995 188.605 ;
        RECT 100.210 188.590 100.530 188.650 ;
        RECT 102.645 188.605 103.295 188.650 ;
        RECT 100.785 188.450 101.075 188.495 ;
        RECT 104.365 188.450 104.655 188.495 ;
        RECT 106.200 188.450 106.490 188.495 ;
        RECT 100.785 188.310 106.490 188.450 ;
        RECT 100.785 188.265 101.075 188.310 ;
        RECT 104.365 188.265 104.655 188.310 ;
        RECT 106.200 188.265 106.490 188.310 ;
        RECT 109.870 188.250 110.190 188.510 ;
        RECT 113.090 188.250 113.410 188.510 ;
        RECT 90.090 188.110 90.410 188.170 ;
        RECT 91.010 188.110 91.330 188.170 ;
        RECT 87.880 187.970 91.330 188.110 ;
        RECT 62.030 187.910 62.350 187.970 ;
        RECT 64.345 187.925 64.635 187.970 ;
        RECT 65.710 187.910 66.030 187.970 ;
        RECT 72.150 187.910 72.470 187.970 ;
        RECT 90.090 187.910 90.410 187.970 ;
        RECT 91.010 187.910 91.330 187.970 ;
        RECT 106.665 188.110 106.955 188.155 ;
        RECT 118.150 188.110 118.470 188.170 ;
        RECT 106.665 187.970 118.470 188.110 ;
        RECT 106.665 187.925 106.955 187.970 ;
        RECT 118.150 187.910 118.470 187.970 ;
        RECT 49.150 187.770 49.470 187.830 ;
        RECT 59.270 187.770 59.590 187.830 ;
        RECT 46.480 187.630 59.590 187.770 ;
        RECT 40.525 187.585 40.815 187.630 ;
        RECT 43.645 187.585 43.935 187.630 ;
        RECT 45.535 187.585 45.825 187.630 ;
        RECT 49.150 187.570 49.470 187.630 ;
        RECT 59.270 187.570 59.590 187.630 ;
        RECT 100.785 187.770 101.075 187.815 ;
        RECT 103.905 187.770 104.195 187.815 ;
        RECT 105.795 187.770 106.085 187.815 ;
        RECT 100.785 187.630 106.085 187.770 ;
        RECT 100.785 187.585 101.075 187.630 ;
        RECT 103.905 187.585 104.195 187.630 ;
        RECT 105.795 187.585 106.085 187.630 ;
        RECT 37.650 187.230 37.970 187.490 ;
        RECT 45.120 187.430 45.410 187.475 ;
        RECT 50.070 187.430 50.390 187.490 ;
        RECT 45.120 187.290 50.390 187.430 ;
        RECT 45.120 187.245 45.410 187.290 ;
        RECT 50.070 187.230 50.390 187.290 ;
        RECT 97.925 187.430 98.215 187.475 ;
        RECT 99.290 187.430 99.610 187.490 ;
        RECT 97.925 187.290 99.610 187.430 ;
        RECT 97.925 187.245 98.215 187.290 ;
        RECT 99.290 187.230 99.610 187.290 ;
        RECT 99.750 187.430 100.070 187.490 ;
        RECT 105.350 187.430 105.640 187.475 ;
        RECT 99.750 187.290 105.640 187.430 ;
        RECT 99.750 187.230 100.070 187.290 ;
        RECT 105.350 187.245 105.640 187.290 ;
        RECT 14.580 186.610 127.740 187.090 ;
        RECT 39.030 186.210 39.350 186.470 ;
        RECT 45.930 186.410 46.250 186.470 ;
        RECT 88.265 186.410 88.555 186.455 ;
        RECT 89.170 186.410 89.490 186.470 ;
        RECT 45.930 186.270 47.540 186.410 ;
        RECT 45.930 186.210 46.250 186.270 ;
        RECT 29.025 186.070 29.315 186.115 ;
        RECT 32.145 186.070 32.435 186.115 ;
        RECT 34.035 186.070 34.325 186.115 ;
        RECT 44.550 186.070 44.870 186.130 ;
        RECT 29.025 185.930 34.325 186.070 ;
        RECT 29.025 185.885 29.315 185.930 ;
        RECT 32.145 185.885 32.435 185.930 ;
        RECT 34.035 185.885 34.325 185.930 ;
        RECT 34.980 185.930 44.870 186.070 ;
        RECT 22.930 185.730 23.250 185.790 ;
        RECT 34.980 185.775 35.120 185.930 ;
        RECT 44.550 185.870 44.870 185.930 ;
        RECT 46.390 185.870 46.710 186.130 ;
        RECT 33.525 185.730 33.815 185.775 ;
        RECT 22.930 185.590 33.815 185.730 ;
        RECT 22.930 185.530 23.250 185.590 ;
        RECT 33.525 185.545 33.815 185.590 ;
        RECT 34.905 185.545 35.195 185.775 ;
        RECT 38.110 185.730 38.430 185.790 ;
        RECT 40.425 185.730 40.715 185.775 ;
        RECT 38.110 185.590 40.715 185.730 ;
        RECT 38.110 185.530 38.430 185.590 ;
        RECT 40.425 185.545 40.715 185.590 ;
        RECT 27.945 185.095 28.235 185.410 ;
        RECT 29.025 185.390 29.315 185.435 ;
        RECT 32.605 185.390 32.895 185.435 ;
        RECT 34.440 185.390 34.730 185.435 ;
        RECT 29.025 185.250 34.730 185.390 ;
        RECT 29.025 185.205 29.315 185.250 ;
        RECT 32.605 185.205 32.895 185.250 ;
        RECT 34.440 185.205 34.730 185.250 ;
        RECT 36.270 185.390 36.590 185.450 ;
        RECT 38.585 185.390 38.875 185.435 ;
        RECT 36.270 185.250 38.875 185.390 ;
        RECT 40.500 185.390 40.640 185.545 ;
        RECT 41.330 185.530 41.650 185.790 ;
        RECT 46.480 185.730 46.620 185.870 ;
        RECT 46.865 185.730 47.155 185.775 ;
        RECT 46.020 185.590 47.155 185.730 ;
        RECT 45.470 185.390 45.790 185.450 ;
        RECT 46.020 185.390 46.160 185.590 ;
        RECT 46.865 185.545 47.155 185.590 ;
        RECT 40.500 185.250 46.160 185.390 ;
        RECT 36.270 185.190 36.590 185.250 ;
        RECT 38.585 185.205 38.875 185.250 ;
        RECT 45.470 185.190 45.790 185.250 ;
        RECT 46.405 185.205 46.695 185.435 ;
        RECT 47.400 185.390 47.540 186.270 ;
        RECT 88.265 186.270 89.490 186.410 ;
        RECT 88.265 186.225 88.555 186.270 ;
        RECT 89.170 186.210 89.490 186.270 ;
        RECT 99.750 186.210 100.070 186.470 ;
        RECT 100.210 186.410 100.530 186.470 ;
        RECT 100.685 186.410 100.975 186.455 ;
        RECT 100.210 186.270 100.975 186.410 ;
        RECT 100.210 186.210 100.530 186.270 ;
        RECT 100.685 186.225 100.975 186.270 ;
        RECT 53.405 186.070 53.695 186.115 ;
        RECT 56.525 186.070 56.815 186.115 ;
        RECT 58.415 186.070 58.705 186.115 ;
        RECT 60.650 186.070 60.970 186.130 ;
        RECT 53.405 185.930 58.705 186.070 ;
        RECT 53.405 185.885 53.695 185.930 ;
        RECT 56.525 185.885 56.815 185.930 ;
        RECT 58.415 185.885 58.705 185.930 ;
        RECT 58.900 185.930 60.970 186.070 ;
        RECT 58.900 185.730 59.040 185.930 ;
        RECT 60.650 185.870 60.970 185.930 ;
        RECT 71.230 186.070 71.550 186.130 ;
        RECT 74.925 186.070 75.215 186.115 ;
        RECT 76.290 186.070 76.610 186.130 ;
        RECT 71.230 185.930 76.610 186.070 ;
        RECT 71.230 185.870 71.550 185.930 ;
        RECT 74.925 185.885 75.215 185.930 ;
        RECT 76.290 185.870 76.610 185.930 ;
        RECT 91.010 186.070 91.330 186.130 ;
        RECT 91.010 185.930 100.440 186.070 ;
        RECT 91.010 185.870 91.330 185.930 ;
        RECT 52.000 185.590 59.040 185.730 ;
        RECT 48.705 185.390 48.995 185.435 ;
        RECT 52.000 185.390 52.140 185.590 ;
        RECT 59.270 185.530 59.590 185.790 ;
        RECT 68.010 185.730 68.330 185.790 ;
        RECT 72.625 185.730 72.915 185.775 ;
        RECT 73.530 185.730 73.850 185.790 ;
        RECT 68.010 185.590 73.850 185.730 ;
        RECT 68.010 185.530 68.330 185.590 ;
        RECT 72.625 185.545 72.915 185.590 ;
        RECT 73.530 185.530 73.850 185.590 ;
        RECT 85.030 185.530 85.350 185.790 ;
        RECT 94.705 185.730 94.995 185.775 ;
        RECT 99.290 185.730 99.610 185.790 ;
        RECT 94.705 185.590 99.610 185.730 ;
        RECT 94.705 185.545 94.995 185.590 ;
        RECT 99.290 185.530 99.610 185.590 ;
        RECT 47.400 185.250 52.140 185.390 ;
        RECT 48.705 185.205 48.995 185.250 ;
        RECT 27.645 185.050 28.235 185.095 ;
        RECT 28.450 185.050 28.770 185.110 ;
        RECT 30.885 185.050 31.535 185.095 ;
        RECT 27.645 184.910 31.535 185.050 ;
        RECT 27.645 184.865 27.935 184.910 ;
        RECT 28.450 184.850 28.770 184.910 ;
        RECT 30.885 184.865 31.535 184.910 ;
        RECT 37.650 185.050 37.970 185.110 ;
        RECT 46.480 185.050 46.620 185.205 ;
        RECT 52.325 185.095 52.615 185.410 ;
        RECT 53.405 185.390 53.695 185.435 ;
        RECT 56.985 185.390 57.275 185.435 ;
        RECT 58.820 185.390 59.110 185.435 ;
        RECT 53.405 185.250 59.110 185.390 ;
        RECT 53.405 185.205 53.695 185.250 ;
        RECT 56.985 185.205 57.275 185.250 ;
        RECT 58.820 185.205 59.110 185.250 ;
        RECT 74.450 185.190 74.770 185.450 ;
        RECT 100.300 185.435 100.440 185.930 ;
        RECT 105.270 185.730 105.590 185.790 ;
        RECT 107.125 185.730 107.415 185.775 ;
        RECT 108.950 185.730 109.270 185.790 ;
        RECT 105.270 185.590 109.270 185.730 ;
        RECT 105.270 185.530 105.590 185.590 ;
        RECT 107.125 185.545 107.415 185.590 ;
        RECT 108.950 185.530 109.270 185.590 ;
        RECT 98.845 185.205 99.135 185.435 ;
        RECT 100.225 185.205 100.515 185.435 ;
        RECT 37.650 184.910 46.620 185.050 ;
        RECT 49.165 185.050 49.455 185.095 ;
        RECT 52.025 185.050 52.615 185.095 ;
        RECT 55.265 185.050 55.915 185.095 ;
        RECT 49.165 184.910 55.915 185.050 ;
        RECT 37.650 184.850 37.970 184.910 ;
        RECT 49.165 184.865 49.455 184.910 ;
        RECT 52.025 184.865 52.315 184.910 ;
        RECT 55.265 184.865 55.915 184.910 ;
        RECT 57.890 184.850 58.210 185.110 ;
        RECT 72.165 185.050 72.455 185.095 ;
        RECT 72.610 185.050 72.930 185.110 ;
        RECT 72.165 184.910 72.930 185.050 ;
        RECT 74.540 185.050 74.680 185.190 ;
        RECT 74.925 185.050 75.215 185.095 ;
        RECT 75.830 185.050 76.150 185.110 ;
        RECT 74.540 184.910 76.150 185.050 ;
        RECT 98.920 185.050 99.060 185.205 ;
        RECT 105.730 185.190 106.050 185.450 ;
        RECT 110.330 185.190 110.650 185.450 ;
        RECT 102.525 185.050 102.815 185.095 ;
        RECT 98.920 184.910 102.815 185.050 ;
        RECT 72.165 184.865 72.455 184.910 ;
        RECT 72.610 184.850 72.930 184.910 ;
        RECT 74.925 184.865 75.215 184.910 ;
        RECT 75.830 184.850 76.150 184.910 ;
        RECT 102.525 184.865 102.815 184.910 ;
        RECT 109.885 185.050 110.175 185.095 ;
        RECT 112.170 185.050 112.490 185.110 ;
        RECT 109.885 184.910 112.490 185.050 ;
        RECT 109.885 184.865 110.175 184.910 ;
        RECT 112.170 184.850 112.490 184.910 ;
        RECT 26.165 184.710 26.455 184.755 ;
        RECT 29.830 184.710 30.150 184.770 ;
        RECT 26.165 184.570 30.150 184.710 ;
        RECT 26.165 184.525 26.455 184.570 ;
        RECT 29.830 184.510 30.150 184.570 ;
        RECT 30.290 184.710 30.610 184.770 ;
        RECT 41.805 184.710 42.095 184.755 ;
        RECT 30.290 184.570 42.095 184.710 ;
        RECT 30.290 184.510 30.610 184.570 ;
        RECT 41.805 184.525 42.095 184.570 ;
        RECT 43.630 184.510 43.950 184.770 ;
        RECT 44.090 184.510 44.410 184.770 ;
        RECT 45.930 184.510 46.250 184.770 ;
        RECT 46.390 184.710 46.710 184.770 ;
        RECT 50.545 184.710 50.835 184.755 ;
        RECT 46.390 184.570 50.835 184.710 ;
        RECT 46.390 184.510 46.710 184.570 ;
        RECT 50.545 184.525 50.835 184.570 ;
        RECT 71.245 184.710 71.535 184.755 ;
        RECT 74.450 184.710 74.770 184.770 ;
        RECT 71.245 184.570 74.770 184.710 ;
        RECT 71.245 184.525 71.535 184.570 ;
        RECT 74.450 184.510 74.770 184.570 ;
        RECT 85.950 184.510 86.270 184.770 ;
        RECT 86.410 184.510 86.730 184.770 ;
        RECT 97.450 184.510 97.770 184.770 ;
        RECT 111.710 184.710 112.030 184.770 ;
        RECT 113.565 184.710 113.855 184.755 ;
        RECT 111.710 184.570 113.855 184.710 ;
        RECT 111.710 184.510 112.030 184.570 ;
        RECT 113.565 184.525 113.855 184.570 ;
        RECT 14.580 183.890 127.740 184.370 ;
        RECT 22.930 183.490 23.250 183.750 ;
        RECT 30.290 183.490 30.610 183.750 ;
        RECT 45.010 183.690 45.330 183.750 ;
        RECT 48.705 183.690 48.995 183.735 ;
        RECT 45.010 183.550 48.995 183.690 ;
        RECT 45.010 183.490 45.330 183.550 ;
        RECT 48.705 183.505 48.995 183.550 ;
        RECT 50.070 183.490 50.390 183.750 ;
        RECT 52.385 183.690 52.675 183.735 ;
        RECT 57.890 183.690 58.210 183.750 ;
        RECT 71.230 183.690 71.550 183.750 ;
        RECT 52.385 183.550 58.210 183.690 ;
        RECT 52.385 183.505 52.675 183.550 ;
        RECT 57.890 183.490 58.210 183.550 ;
        RECT 69.020 183.550 71.550 183.690 ;
        RECT 32.605 183.350 32.895 183.395 ;
        RECT 33.970 183.350 34.290 183.410 ;
        RECT 32.605 183.210 34.290 183.350 ;
        RECT 32.605 183.165 32.895 183.210 ;
        RECT 33.970 183.150 34.290 183.210 ;
        RECT 44.565 183.350 44.855 183.395 ;
        RECT 44.565 183.210 51.220 183.350 ;
        RECT 44.565 183.165 44.855 183.210 ;
        RECT 22.025 183.010 22.315 183.055 ;
        RECT 23.405 183.010 23.695 183.055 ;
        RECT 22.025 182.870 23.695 183.010 ;
        RECT 22.025 182.825 22.315 182.870 ;
        RECT 23.405 182.825 23.695 182.870 ;
        RECT 27.545 183.010 27.835 183.055 ;
        RECT 29.830 183.010 30.150 183.070 ;
        RECT 33.065 183.010 33.355 183.055 ;
        RECT 35.810 183.010 36.130 183.070 ;
        RECT 27.545 182.870 36.130 183.010 ;
        RECT 27.545 182.825 27.835 182.870 ;
        RECT 29.830 182.810 30.150 182.870 ;
        RECT 33.065 182.825 33.355 182.870 ;
        RECT 35.810 182.810 36.130 182.870 ;
        RECT 37.650 182.810 37.970 183.070 ;
        RECT 41.805 183.010 42.095 183.055 ;
        RECT 44.090 183.010 44.410 183.070 ;
        RECT 41.805 182.870 44.410 183.010 ;
        RECT 41.805 182.825 42.095 182.870 ;
        RECT 44.090 182.810 44.410 182.870 ;
        RECT 45.485 183.010 45.775 183.055 ;
        RECT 46.390 183.010 46.710 183.070 ;
        RECT 51.080 183.055 51.220 183.210 ;
        RECT 45.485 182.870 46.710 183.010 ;
        RECT 45.485 182.825 45.775 182.870 ;
        RECT 46.390 182.810 46.710 182.870 ;
        RECT 49.625 182.825 49.915 183.055 ;
        RECT 51.005 182.825 51.295 183.055 ;
        RECT 51.465 182.825 51.755 183.055 ;
        RECT 55.605 183.010 55.895 183.055 ;
        RECT 59.270 183.010 59.590 183.070 ;
        RECT 55.605 182.870 59.590 183.010 ;
        RECT 55.605 182.825 55.895 182.870 ;
        RECT 26.625 182.485 26.915 182.715 ;
        RECT 33.985 182.670 34.275 182.715 ;
        RECT 38.110 182.670 38.430 182.730 ;
        RECT 33.985 182.530 38.430 182.670 ;
        RECT 33.985 182.485 34.275 182.530 ;
        RECT 26.700 182.330 26.840 182.485 ;
        RECT 38.110 182.470 38.430 182.530 ;
        RECT 43.630 182.670 43.950 182.730 ;
        RECT 49.700 182.670 49.840 182.825 ;
        RECT 43.630 182.530 49.840 182.670 ;
        RECT 50.070 182.670 50.390 182.730 ;
        RECT 51.540 182.670 51.680 182.825 ;
        RECT 59.270 182.810 59.590 182.870 ;
        RECT 60.205 183.010 60.495 183.055 ;
        RECT 60.650 183.010 60.970 183.070 ;
        RECT 60.205 182.870 60.970 183.010 ;
        RECT 60.205 182.825 60.495 182.870 ;
        RECT 60.650 182.810 60.970 182.870 ;
        RECT 68.010 182.810 68.330 183.070 ;
        RECT 69.020 183.055 69.160 183.550 ;
        RECT 71.230 183.490 71.550 183.550 ;
        RECT 71.690 183.690 72.010 183.750 ;
        RECT 72.610 183.690 72.930 183.750 ;
        RECT 73.990 183.690 74.310 183.750 ;
        RECT 89.645 183.690 89.935 183.735 ;
        RECT 71.690 183.550 76.520 183.690 ;
        RECT 71.690 183.490 72.010 183.550 ;
        RECT 72.610 183.490 72.930 183.550 ;
        RECT 73.990 183.490 74.310 183.550 ;
        RECT 73.530 183.150 73.850 183.410 ;
        RECT 68.945 182.825 69.235 183.055 ;
        RECT 70.785 183.010 71.075 183.055 ;
        RECT 71.690 183.010 72.010 183.070 ;
        RECT 70.785 182.870 72.010 183.010 ;
        RECT 70.785 182.825 71.075 182.870 ;
        RECT 50.070 182.530 51.680 182.670 ;
        RECT 43.630 182.470 43.950 182.530 ;
        RECT 50.070 182.470 50.390 182.530 ;
        RECT 67.565 182.485 67.855 182.715 ;
        RECT 68.485 182.670 68.775 182.715 ;
        RECT 70.860 182.670 71.000 182.825 ;
        RECT 71.690 182.810 72.010 182.870 ;
        RECT 72.165 182.825 72.455 183.055 ;
        RECT 68.485 182.530 71.000 182.670 ;
        RECT 72.240 182.670 72.380 182.825 ;
        RECT 72.610 182.810 72.930 183.070 ;
        RECT 73.620 183.010 73.760 183.150 ;
        RECT 74.925 183.010 75.215 183.055 ;
        RECT 73.620 182.870 75.215 183.010 ;
        RECT 74.925 182.825 75.215 182.870 ;
        RECT 72.240 182.530 72.840 182.670 ;
        RECT 68.485 182.485 68.775 182.530 ;
        RECT 30.765 182.330 31.055 182.375 ;
        RECT 26.700 182.190 31.055 182.330 ;
        RECT 67.640 182.330 67.780 182.485 ;
        RECT 72.700 182.390 72.840 182.530 ;
        RECT 73.530 182.470 73.850 182.730 ;
        RECT 75.000 182.670 75.140 182.825 ;
        RECT 75.830 182.810 76.150 183.070 ;
        RECT 76.380 183.055 76.520 183.550 ;
        RECT 86.500 183.550 89.935 183.690 ;
        RECT 81.005 183.350 81.295 183.395 ;
        RECT 84.245 183.350 84.895 183.395 ;
        RECT 86.500 183.350 86.640 183.550 ;
        RECT 89.645 183.505 89.935 183.550 ;
        RECT 97.450 183.490 97.770 183.750 ;
        RECT 105.730 183.690 106.050 183.750 ;
        RECT 106.205 183.690 106.495 183.735 ;
        RECT 105.730 183.550 106.495 183.690 ;
        RECT 105.730 183.490 106.050 183.550 ;
        RECT 106.205 183.505 106.495 183.550 ;
        RECT 111.725 183.505 112.015 183.735 ;
        RECT 81.005 183.210 86.640 183.350 ;
        RECT 104.365 183.350 104.655 183.395 ;
        RECT 111.800 183.350 111.940 183.505 ;
        RECT 104.365 183.210 111.940 183.350 ;
        RECT 117.345 183.350 117.635 183.395 ;
        RECT 120.585 183.350 121.235 183.395 ;
        RECT 117.345 183.210 121.235 183.350 ;
        RECT 81.005 183.165 81.595 183.210 ;
        RECT 84.245 183.165 84.895 183.210 ;
        RECT 104.365 183.165 104.655 183.210 ;
        RECT 76.305 182.825 76.595 183.055 ;
        RECT 76.750 182.810 77.070 183.070 ;
        RECT 81.305 182.850 81.595 183.165 ;
        RECT 105.820 183.070 105.960 183.210 ;
        RECT 117.345 183.165 117.935 183.210 ;
        RECT 120.585 183.165 121.235 183.210 ;
        RECT 123.225 183.350 123.515 183.395 ;
        RECT 124.590 183.350 124.910 183.410 ;
        RECT 123.225 183.210 124.910 183.350 ;
        RECT 123.225 183.165 123.515 183.210 ;
        RECT 117.645 183.070 117.935 183.165 ;
        RECT 124.590 183.150 124.910 183.210 ;
        RECT 82.385 183.010 82.675 183.055 ;
        RECT 85.965 183.010 86.255 183.055 ;
        RECT 87.800 183.010 88.090 183.055 ;
        RECT 82.385 182.870 88.090 183.010 ;
        RECT 82.385 182.825 82.675 182.870 ;
        RECT 85.965 182.825 86.255 182.870 ;
        RECT 87.800 182.825 88.090 182.870 ;
        RECT 90.105 183.010 90.395 183.055 ;
        RECT 91.010 183.010 91.330 183.070 ;
        RECT 90.105 182.870 91.330 183.010 ;
        RECT 90.105 182.825 90.395 182.870 ;
        RECT 91.010 182.810 91.330 182.870 ;
        RECT 96.070 183.010 96.390 183.070 ;
        RECT 97.005 183.010 97.295 183.055 ;
        RECT 96.070 182.870 97.295 183.010 ;
        RECT 96.070 182.810 96.390 182.870 ;
        RECT 97.005 182.825 97.295 182.870 ;
        RECT 99.290 183.010 99.610 183.070 ;
        RECT 103.905 183.010 104.195 183.055 ;
        RECT 99.290 182.870 104.195 183.010 ;
        RECT 99.290 182.810 99.610 182.870 ;
        RECT 103.905 182.825 104.195 182.870 ;
        RECT 105.730 182.810 106.050 183.070 ;
        RECT 106.190 183.010 106.510 183.070 ;
        RECT 106.190 182.870 107.800 183.010 ;
        RECT 106.190 182.810 106.510 182.870 ;
        RECT 77.225 182.670 77.515 182.715 ;
        RECT 75.000 182.530 77.515 182.670 ;
        RECT 77.225 182.485 77.515 182.530 ;
        RECT 86.885 182.670 87.175 182.715 ;
        RECT 88.265 182.670 88.555 182.715 ;
        RECT 93.770 182.670 94.090 182.730 ;
        RECT 86.885 182.530 88.020 182.670 ;
        RECT 86.885 182.485 87.175 182.530 ;
        RECT 72.610 182.330 72.930 182.390 ;
        RECT 75.830 182.330 76.150 182.390 ;
        RECT 67.640 182.190 76.150 182.330 ;
        RECT 30.765 182.145 31.055 182.190 ;
        RECT 72.610 182.130 72.930 182.190 ;
        RECT 75.830 182.130 76.150 182.190 ;
        RECT 82.385 182.330 82.675 182.375 ;
        RECT 85.505 182.330 85.795 182.375 ;
        RECT 87.395 182.330 87.685 182.375 ;
        RECT 82.385 182.190 87.685 182.330 ;
        RECT 87.880 182.330 88.020 182.530 ;
        RECT 88.265 182.530 94.090 182.670 ;
        RECT 88.265 182.485 88.555 182.530 ;
        RECT 93.770 182.470 94.090 182.530 ;
        RECT 96.545 182.670 96.835 182.715 ;
        RECT 97.910 182.670 98.230 182.730 ;
        RECT 102.985 182.670 103.275 182.715 ;
        RECT 96.545 182.530 103.275 182.670 ;
        RECT 96.545 182.485 96.835 182.530 ;
        RECT 89.630 182.330 89.950 182.390 ;
        RECT 87.880 182.190 89.950 182.330 ;
        RECT 82.385 182.145 82.675 182.190 ;
        RECT 85.505 182.145 85.795 182.190 ;
        RECT 87.395 182.145 87.685 182.190 ;
        RECT 89.630 182.130 89.950 182.190 ;
        RECT 39.490 181.990 39.810 182.050 ;
        RECT 40.885 181.990 41.175 182.035 ;
        RECT 39.490 181.850 41.175 181.990 ;
        RECT 39.490 181.790 39.810 181.850 ;
        RECT 40.885 181.805 41.175 181.850 ;
        RECT 45.930 181.990 46.250 182.050 ;
        RECT 47.310 181.990 47.630 182.050 ;
        RECT 48.245 181.990 48.535 182.035 ;
        RECT 45.930 181.850 48.535 181.990 ;
        RECT 45.930 181.790 46.250 181.850 ;
        RECT 47.310 181.790 47.630 181.850 ;
        RECT 48.245 181.805 48.535 181.850 ;
        RECT 56.050 181.990 56.370 182.050 ;
        RECT 59.745 181.990 60.035 182.035 ;
        RECT 56.050 181.850 60.035 181.990 ;
        RECT 56.050 181.790 56.370 181.850 ;
        RECT 59.745 181.805 60.035 181.850 ;
        RECT 66.645 181.990 66.935 182.035 ;
        RECT 69.390 181.990 69.710 182.050 ;
        RECT 66.645 181.850 69.710 181.990 ;
        RECT 66.645 181.805 66.935 181.850 ;
        RECT 69.390 181.790 69.710 181.850 ;
        RECT 74.910 181.990 75.230 182.050 ;
        RECT 78.145 181.990 78.435 182.035 ;
        RECT 74.910 181.850 78.435 181.990 ;
        RECT 74.910 181.790 75.230 181.850 ;
        RECT 78.145 181.805 78.435 181.850 ;
        RECT 79.510 181.790 79.830 182.050 ;
        RECT 85.030 181.990 85.350 182.050 ;
        RECT 96.620 181.990 96.760 182.485 ;
        RECT 97.910 182.470 98.230 182.530 ;
        RECT 102.985 182.485 103.275 182.530 ;
        RECT 104.350 182.670 104.670 182.730 ;
        RECT 106.665 182.670 106.955 182.715 ;
        RECT 104.350 182.530 106.955 182.670 ;
        RECT 107.660 182.670 107.800 182.870 ;
        RECT 108.030 182.810 108.350 183.070 ;
        RECT 108.505 182.825 108.795 183.055 ;
        RECT 108.965 182.825 109.255 183.055 ;
        RECT 109.410 183.010 109.730 183.070 ;
        RECT 109.885 183.010 110.175 183.055 ;
        RECT 109.410 182.870 110.175 183.010 ;
        RECT 108.580 182.670 108.720 182.825 ;
        RECT 107.660 182.530 108.720 182.670 ;
        RECT 104.350 182.470 104.670 182.530 ;
        RECT 106.665 182.485 106.955 182.530 ;
        RECT 98.370 182.330 98.690 182.390 ;
        RECT 109.040 182.330 109.180 182.825 ;
        RECT 109.410 182.810 109.730 182.870 ;
        RECT 109.885 182.825 110.175 182.870 ;
        RECT 111.710 183.010 112.030 183.070 ;
        RECT 112.185 183.010 112.475 183.055 ;
        RECT 111.710 182.870 112.475 183.010 ;
        RECT 111.710 182.810 112.030 182.870 ;
        RECT 112.185 182.825 112.475 182.870 ;
        RECT 117.645 182.850 118.010 183.070 ;
        RECT 117.690 182.810 118.010 182.850 ;
        RECT 118.725 183.010 119.015 183.055 ;
        RECT 122.305 183.010 122.595 183.055 ;
        RECT 124.140 183.010 124.430 183.055 ;
        RECT 118.725 182.870 124.430 183.010 ;
        RECT 118.725 182.825 119.015 182.870 ;
        RECT 122.305 182.825 122.595 182.870 ;
        RECT 124.140 182.825 124.430 182.870 ;
        RECT 110.790 182.470 111.110 182.730 ;
        RECT 118.150 182.670 118.470 182.730 ;
        RECT 124.605 182.670 124.895 182.715 ;
        RECT 118.150 182.530 124.895 182.670 ;
        RECT 118.150 182.470 118.470 182.530 ;
        RECT 124.605 182.485 124.895 182.530 ;
        RECT 98.370 182.190 109.180 182.330 ;
        RECT 110.330 182.330 110.650 182.390 ;
        RECT 115.865 182.330 116.155 182.375 ;
        RECT 110.330 182.190 116.155 182.330 ;
        RECT 98.370 182.130 98.690 182.190 ;
        RECT 110.330 182.130 110.650 182.190 ;
        RECT 115.865 182.145 116.155 182.190 ;
        RECT 118.725 182.330 119.015 182.375 ;
        RECT 121.845 182.330 122.135 182.375 ;
        RECT 123.735 182.330 124.025 182.375 ;
        RECT 118.725 182.190 124.025 182.330 ;
        RECT 118.725 182.145 119.015 182.190 ;
        RECT 121.845 182.145 122.135 182.190 ;
        RECT 123.735 182.145 124.025 182.190 ;
        RECT 85.030 181.850 96.760 181.990 ;
        RECT 99.305 181.990 99.595 182.035 ;
        RECT 104.810 181.990 105.130 182.050 ;
        RECT 99.305 181.850 105.130 181.990 ;
        RECT 85.030 181.790 85.350 181.850 ;
        RECT 99.305 181.805 99.595 181.850 ;
        RECT 104.810 181.790 105.130 181.850 ;
        RECT 114.025 181.990 114.315 182.035 ;
        RECT 116.770 181.990 117.090 182.050 ;
        RECT 114.025 181.850 117.090 181.990 ;
        RECT 114.025 181.805 114.315 181.850 ;
        RECT 116.770 181.790 117.090 181.850 ;
        RECT 14.580 181.170 127.740 181.650 ;
        RECT 45.470 180.970 45.790 181.030 ;
        RECT 46.850 180.970 47.170 181.030 ;
        RECT 45.470 180.830 47.170 180.970 ;
        RECT 45.470 180.770 45.790 180.830 ;
        RECT 46.850 180.770 47.170 180.830 ;
        RECT 49.625 180.970 49.915 181.015 ;
        RECT 50.070 180.970 50.390 181.030 ;
        RECT 82.270 180.970 82.590 181.030 ;
        RECT 49.625 180.830 50.390 180.970 ;
        RECT 49.625 180.785 49.915 180.830 ;
        RECT 50.070 180.770 50.390 180.830 ;
        RECT 78.680 180.830 82.590 180.970 ;
        RECT 25.655 180.630 25.945 180.675 ;
        RECT 27.545 180.630 27.835 180.675 ;
        RECT 30.665 180.630 30.955 180.675 ;
        RECT 25.655 180.490 30.955 180.630 ;
        RECT 25.655 180.445 25.945 180.490 ;
        RECT 27.545 180.445 27.835 180.490 ;
        RECT 30.665 180.445 30.955 180.490 ;
        RECT 53.765 180.630 54.055 180.675 ;
        RECT 56.510 180.630 56.830 180.690 ;
        RECT 53.765 180.490 56.830 180.630 ;
        RECT 53.765 180.445 54.055 180.490 ;
        RECT 56.510 180.430 56.830 180.490 ;
        RECT 67.550 180.630 67.870 180.690 ;
        RECT 78.680 180.630 78.820 180.830 ;
        RECT 82.270 180.770 82.590 180.830 ;
        RECT 89.630 180.770 89.950 181.030 ;
        RECT 105.730 180.770 106.050 181.030 ;
        RECT 117.690 180.970 118.010 181.030 ;
        RECT 122.765 180.970 123.055 181.015 ;
        RECT 124.590 180.970 124.910 181.030 ;
        RECT 117.690 180.830 119.760 180.970 ;
        RECT 117.690 180.770 118.010 180.830 ;
        RECT 67.550 180.490 78.820 180.630 ;
        RECT 79.050 180.630 79.370 180.690 ;
        RECT 85.490 180.630 85.810 180.690 ;
        RECT 79.050 180.490 85.810 180.630 ;
        RECT 67.550 180.430 67.870 180.490 ;
        RECT 79.050 180.430 79.370 180.490 ;
        RECT 85.490 180.430 85.810 180.490 ;
        RECT 95.265 180.630 95.555 180.675 ;
        RECT 98.385 180.630 98.675 180.675 ;
        RECT 100.275 180.630 100.565 180.675 ;
        RECT 95.265 180.490 100.565 180.630 ;
        RECT 95.265 180.445 95.555 180.490 ;
        RECT 98.385 180.445 98.675 180.490 ;
        RECT 100.275 180.445 100.565 180.490 ;
        RECT 114.125 180.630 114.415 180.675 ;
        RECT 117.245 180.630 117.535 180.675 ;
        RECT 119.135 180.630 119.425 180.675 ;
        RECT 114.125 180.490 119.425 180.630 ;
        RECT 119.620 180.630 119.760 180.830 ;
        RECT 122.765 180.830 124.910 180.970 ;
        RECT 122.765 180.785 123.055 180.830 ;
        RECT 124.590 180.770 124.910 180.830 ;
        RECT 120.925 180.630 121.215 180.675 ;
        RECT 119.620 180.490 121.215 180.630 ;
        RECT 114.125 180.445 114.415 180.490 ;
        RECT 117.245 180.445 117.535 180.490 ;
        RECT 119.135 180.445 119.425 180.490 ;
        RECT 120.925 180.445 121.215 180.490 ;
        RECT 33.525 180.105 33.815 180.335 ;
        RECT 46.390 180.290 46.710 180.350 ;
        RECT 44.640 180.150 46.710 180.290 ;
        RECT 24.785 179.765 25.075 179.995 ;
        RECT 25.250 179.950 25.540 179.995 ;
        RECT 27.085 179.950 27.375 179.995 ;
        RECT 30.665 179.950 30.955 179.995 ;
        RECT 25.250 179.810 30.955 179.950 ;
        RECT 25.250 179.765 25.540 179.810 ;
        RECT 27.085 179.765 27.375 179.810 ;
        RECT 30.665 179.765 30.955 179.810 ;
        RECT 24.860 179.610 25.000 179.765 ;
        RECT 24.860 179.470 25.460 179.610 ;
        RECT 25.320 179.270 25.460 179.470 ;
        RECT 26.150 179.410 26.470 179.670 ;
        RECT 27.530 179.610 27.850 179.670 ;
        RECT 31.745 179.655 32.035 179.970 ;
        RECT 33.600 179.950 33.740 180.105 ;
        RECT 37.190 179.950 37.510 180.010 ;
        RECT 33.600 179.810 37.510 179.950 ;
        RECT 37.190 179.750 37.510 179.810 ;
        RECT 39.505 179.765 39.795 179.995 ;
        RECT 39.965 179.765 40.255 179.995 ;
        RECT 40.425 179.950 40.715 179.995 ;
        RECT 40.870 179.950 41.190 180.010 ;
        RECT 40.425 179.810 41.190 179.950 ;
        RECT 40.425 179.765 40.715 179.810 ;
        RECT 28.445 179.610 29.095 179.655 ;
        RECT 31.745 179.610 32.335 179.655 ;
        RECT 27.530 179.470 32.335 179.610 ;
        RECT 27.530 179.410 27.850 179.470 ;
        RECT 28.445 179.425 29.095 179.470 ;
        RECT 32.045 179.425 32.335 179.470 ;
        RECT 33.970 179.410 34.290 179.670 ;
        RECT 34.890 179.610 35.210 179.670 ;
        RECT 38.125 179.610 38.415 179.655 ;
        RECT 34.890 179.470 38.415 179.610 ;
        RECT 34.890 179.410 35.210 179.470 ;
        RECT 38.125 179.425 38.415 179.470 ;
        RECT 36.730 179.270 37.050 179.330 ;
        RECT 25.320 179.130 37.050 179.270 ;
        RECT 39.580 179.270 39.720 179.765 ;
        RECT 40.040 179.610 40.180 179.765 ;
        RECT 40.870 179.750 41.190 179.810 ;
        RECT 41.345 179.765 41.635 179.995 ;
        RECT 43.645 179.765 43.935 179.995 ;
        RECT 40.040 179.470 40.640 179.610 ;
        RECT 40.500 179.330 40.640 179.470 ;
        RECT 39.950 179.270 40.270 179.330 ;
        RECT 39.580 179.130 40.270 179.270 ;
        RECT 36.730 179.070 37.050 179.130 ;
        RECT 39.950 179.070 40.270 179.130 ;
        RECT 40.410 179.070 40.730 179.330 ;
        RECT 40.870 179.270 41.190 179.330 ;
        RECT 41.420 179.270 41.560 179.765 ;
        RECT 40.870 179.130 41.560 179.270 ;
        RECT 40.870 179.070 41.190 179.130 ;
        RECT 42.250 179.070 42.570 179.330 ;
        RECT 43.720 179.270 43.860 179.765 ;
        RECT 44.090 179.750 44.410 180.010 ;
        RECT 44.640 179.995 44.780 180.150 ;
        RECT 46.390 180.090 46.710 180.150 ;
        RECT 46.850 180.090 47.170 180.350 ;
        RECT 47.310 180.090 47.630 180.350 ;
        RECT 51.005 180.290 51.295 180.335 ;
        RECT 52.370 180.290 52.690 180.350 ;
        RECT 51.005 180.150 52.690 180.290 ;
        RECT 51.005 180.105 51.295 180.150 ;
        RECT 52.370 180.090 52.690 180.150 ;
        RECT 54.210 180.290 54.530 180.350 ;
        RECT 58.825 180.290 59.115 180.335 ;
        RECT 60.665 180.290 60.955 180.335 ;
        RECT 54.210 180.150 60.955 180.290 ;
        RECT 54.210 180.090 54.530 180.150 ;
        RECT 58.825 180.105 59.115 180.150 ;
        RECT 60.665 180.105 60.955 180.150 ;
        RECT 72.610 180.090 72.930 180.350 ;
        RECT 73.070 180.090 73.390 180.350 ;
        RECT 73.545 180.290 73.835 180.335 ;
        RECT 75.830 180.290 76.150 180.350 ;
        RECT 73.545 180.150 76.150 180.290 ;
        RECT 73.545 180.105 73.835 180.150 ;
        RECT 75.830 180.090 76.150 180.150 ;
        RECT 76.765 180.290 77.055 180.335 ;
        RECT 79.510 180.290 79.830 180.350 ;
        RECT 85.030 180.290 85.350 180.350 ;
        RECT 85.965 180.290 86.255 180.335 ;
        RECT 76.765 180.150 81.120 180.290 ;
        RECT 76.765 180.105 77.055 180.150 ;
        RECT 79.510 180.090 79.830 180.150 ;
        RECT 44.565 179.765 44.855 179.995 ;
        RECT 45.470 179.750 45.790 180.010 ;
        RECT 65.710 179.750 66.030 180.010 ;
        RECT 68.470 179.750 68.790 180.010 ;
        RECT 71.230 179.950 71.550 180.010 ;
        RECT 71.705 179.950 71.995 179.995 ;
        RECT 71.230 179.810 71.995 179.950 ;
        RECT 71.230 179.750 71.550 179.810 ;
        RECT 71.705 179.765 71.995 179.810 ;
        RECT 73.990 179.750 74.310 180.010 ;
        RECT 76.290 179.950 76.610 180.010 ;
        RECT 80.980 179.995 81.120 180.150 ;
        RECT 85.030 180.150 86.255 180.290 ;
        RECT 85.030 180.090 85.350 180.150 ;
        RECT 85.965 180.105 86.255 180.150 ;
        RECT 104.810 180.090 105.130 180.350 ;
        RECT 105.730 180.290 106.050 180.350 ;
        RECT 108.030 180.290 108.350 180.350 ;
        RECT 111.265 180.290 111.555 180.335 ;
        RECT 115.850 180.290 116.170 180.350 ;
        RECT 105.730 180.150 108.350 180.290 ;
        RECT 105.730 180.090 106.050 180.150 ;
        RECT 108.030 180.090 108.350 180.150 ;
        RECT 109.040 180.150 111.555 180.290 ;
        RECT 109.040 180.010 109.180 180.150 ;
        RECT 111.265 180.105 111.555 180.150 ;
        RECT 111.800 180.150 120.680 180.290 ;
        RECT 79.985 179.950 80.275 179.995 ;
        RECT 76.290 179.810 80.275 179.950 ;
        RECT 76.290 179.750 76.610 179.810 ;
        RECT 53.750 179.610 54.070 179.670 ;
        RECT 58.365 179.610 58.655 179.655 ;
        RECT 53.750 179.470 58.655 179.610 ;
        RECT 53.750 179.410 54.070 179.470 ;
        RECT 58.365 179.425 58.655 179.470 ;
        RECT 62.045 179.610 62.335 179.655 ;
        RECT 69.405 179.610 69.695 179.655 ;
        RECT 73.070 179.610 73.390 179.670 ;
        RECT 62.045 179.470 73.390 179.610 ;
        RECT 62.045 179.425 62.335 179.470 ;
        RECT 69.405 179.425 69.695 179.470 ;
        RECT 73.070 179.410 73.390 179.470 ;
        RECT 44.550 179.270 44.870 179.330 ;
        RECT 43.720 179.130 44.870 179.270 ;
        RECT 44.550 179.070 44.870 179.130 ;
        RECT 45.930 179.270 46.250 179.330 ;
        RECT 47.785 179.270 48.075 179.315 ;
        RECT 45.930 179.130 48.075 179.270 ;
        RECT 45.930 179.070 46.250 179.130 ;
        RECT 47.785 179.085 48.075 179.130 ;
        RECT 50.530 179.270 50.850 179.330 ;
        RECT 56.065 179.270 56.355 179.315 ;
        RECT 50.530 179.130 56.355 179.270 ;
        RECT 50.530 179.070 50.850 179.130 ;
        RECT 56.065 179.085 56.355 179.130 ;
        RECT 57.890 179.070 58.210 179.330 ;
        RECT 66.170 179.070 66.490 179.330 ;
        RECT 70.785 179.270 71.075 179.315 ;
        RECT 78.590 179.270 78.910 179.330 ;
        RECT 70.785 179.130 78.910 179.270 ;
        RECT 79.140 179.270 79.280 179.810 ;
        RECT 79.985 179.765 80.275 179.810 ;
        RECT 80.905 179.765 81.195 179.995 ;
        RECT 81.350 179.750 81.670 180.010 ;
        RECT 81.810 179.750 82.130 180.010 ;
        RECT 90.550 179.750 90.870 180.010 ;
        RECT 91.010 179.750 91.330 180.010 ;
        RECT 79.525 179.610 79.815 179.655 ;
        RECT 86.410 179.610 86.730 179.670 ;
        RECT 94.185 179.655 94.475 179.970 ;
        RECT 95.265 179.950 95.555 179.995 ;
        RECT 98.845 179.950 99.135 179.995 ;
        RECT 100.680 179.950 100.970 179.995 ;
        RECT 95.265 179.810 100.970 179.950 ;
        RECT 95.265 179.765 95.555 179.810 ;
        RECT 98.845 179.765 99.135 179.810 ;
        RECT 100.680 179.765 100.970 179.810 ;
        RECT 101.145 179.765 101.435 179.995 ;
        RECT 86.885 179.610 87.175 179.655 ;
        RECT 91.485 179.610 91.775 179.655 ;
        RECT 93.885 179.610 94.475 179.655 ;
        RECT 97.125 179.610 97.775 179.655 ;
        RECT 79.525 179.470 87.175 179.610 ;
        RECT 79.525 179.425 79.815 179.470 ;
        RECT 86.410 179.410 86.730 179.470 ;
        RECT 86.885 179.425 87.175 179.470 ;
        RECT 87.420 179.470 90.320 179.610 ;
        RECT 87.420 179.330 87.560 179.470 ;
        RECT 82.730 179.270 83.050 179.330 ;
        RECT 79.140 179.130 83.050 179.270 ;
        RECT 70.785 179.085 71.075 179.130 ;
        RECT 78.590 179.070 78.910 179.130 ;
        RECT 82.730 179.070 83.050 179.130 ;
        RECT 83.205 179.270 83.495 179.315 ;
        RECT 83.650 179.270 83.970 179.330 ;
        RECT 83.205 179.130 83.970 179.270 ;
        RECT 83.205 179.085 83.495 179.130 ;
        RECT 83.650 179.070 83.970 179.130 ;
        RECT 87.330 179.070 87.650 179.330 ;
        RECT 89.170 179.070 89.490 179.330 ;
        RECT 90.180 179.270 90.320 179.470 ;
        RECT 91.485 179.470 97.775 179.610 ;
        RECT 91.485 179.425 91.775 179.470 ;
        RECT 93.885 179.425 94.175 179.470 ;
        RECT 97.125 179.425 97.775 179.470 ;
        RECT 99.750 179.410 100.070 179.670 ;
        RECT 92.405 179.270 92.695 179.315 ;
        RECT 96.070 179.270 96.390 179.330 ;
        RECT 90.180 179.130 96.390 179.270 ;
        RECT 101.220 179.270 101.360 179.765 ;
        RECT 108.950 179.750 109.270 180.010 ;
        RECT 109.885 179.950 110.175 179.995 ;
        RECT 111.800 179.950 111.940 180.150 ;
        RECT 115.850 180.090 116.170 180.150 ;
        RECT 120.540 179.995 120.680 180.150 ;
        RECT 109.885 179.810 111.940 179.950 ;
        RECT 109.885 179.765 110.175 179.810 ;
        RECT 102.050 179.410 102.370 179.670 ;
        RECT 113.045 179.655 113.335 179.970 ;
        RECT 114.125 179.950 114.415 179.995 ;
        RECT 117.705 179.950 117.995 179.995 ;
        RECT 119.540 179.950 119.830 179.995 ;
        RECT 114.125 179.810 119.830 179.950 ;
        RECT 114.125 179.765 114.415 179.810 ;
        RECT 117.705 179.765 117.995 179.810 ;
        RECT 119.540 179.765 119.830 179.810 ;
        RECT 120.005 179.765 120.295 179.995 ;
        RECT 120.465 179.765 120.755 179.995 ;
        RECT 110.345 179.610 110.635 179.655 ;
        RECT 112.745 179.610 113.335 179.655 ;
        RECT 115.985 179.610 116.635 179.655 ;
        RECT 110.345 179.470 116.635 179.610 ;
        RECT 110.345 179.425 110.635 179.470 ;
        RECT 112.745 179.425 113.035 179.470 ;
        RECT 115.985 179.425 116.635 179.470 ;
        RECT 118.610 179.410 118.930 179.670 ;
        RECT 118.150 179.270 118.470 179.330 ;
        RECT 120.080 179.270 120.220 179.765 ;
        RECT 121.830 179.750 122.150 180.010 ;
        RECT 101.220 179.130 120.220 179.270 ;
        RECT 92.405 179.085 92.695 179.130 ;
        RECT 96.070 179.070 96.390 179.130 ;
        RECT 118.150 179.070 118.470 179.130 ;
        RECT 14.580 178.450 127.740 178.930 ;
        RECT 25.705 178.250 25.995 178.295 ;
        RECT 27.530 178.250 27.850 178.310 ;
        RECT 25.705 178.110 27.850 178.250 ;
        RECT 25.705 178.065 25.995 178.110 ;
        RECT 27.530 178.050 27.850 178.110 ;
        RECT 39.490 178.050 39.810 178.310 ;
        RECT 45.930 178.050 46.250 178.310 ;
        RECT 53.750 178.250 54.070 178.310 ;
        RECT 62.030 178.250 62.350 178.310 ;
        RECT 63.425 178.250 63.715 178.295 ;
        RECT 71.690 178.250 72.010 178.310 ;
        RECT 72.165 178.250 72.455 178.295 ;
        RECT 46.480 178.110 54.070 178.250 ;
        RECT 27.085 177.910 27.375 177.955 ;
        RECT 29.485 177.910 29.775 177.955 ;
        RECT 32.725 177.910 33.375 177.955 ;
        RECT 46.480 177.910 46.620 178.110 ;
        RECT 53.750 178.050 54.070 178.110 ;
        RECT 54.760 178.110 61.800 178.250 ;
        RECT 52.370 177.910 52.690 177.970 ;
        RECT 27.085 177.770 33.375 177.910 ;
        RECT 27.085 177.725 27.375 177.770 ;
        RECT 29.485 177.725 30.075 177.770 ;
        RECT 32.725 177.725 33.375 177.770 ;
        RECT 43.260 177.770 46.620 177.910 ;
        RECT 47.400 177.770 52.690 177.910 ;
        RECT 26.165 177.570 26.455 177.615 ;
        RECT 26.625 177.570 26.915 177.615 ;
        RECT 26.165 177.430 26.915 177.570 ;
        RECT 26.165 177.385 26.455 177.430 ;
        RECT 26.625 177.385 26.915 177.430 ;
        RECT 29.785 177.410 30.075 177.725 ;
        RECT 43.260 177.615 43.400 177.770 ;
        RECT 30.865 177.570 31.155 177.615 ;
        RECT 34.445 177.570 34.735 177.615 ;
        RECT 36.280 177.570 36.570 177.615 ;
        RECT 30.865 177.430 36.570 177.570 ;
        RECT 30.865 177.385 31.155 177.430 ;
        RECT 34.445 177.385 34.735 177.430 ;
        RECT 36.280 177.385 36.570 177.430 ;
        RECT 43.185 177.570 43.475 177.615 ;
        RECT 43.630 177.570 43.950 177.630 ;
        RECT 43.185 177.430 43.950 177.570 ;
        RECT 43.185 177.385 43.475 177.430 ;
        RECT 26.700 177.230 26.840 177.385 ;
        RECT 43.630 177.370 43.950 177.430 ;
        RECT 45.470 177.570 45.790 177.630 ;
        RECT 47.400 177.615 47.540 177.770 ;
        RECT 52.370 177.710 52.690 177.770 ;
        RECT 46.405 177.570 46.695 177.615 ;
        RECT 45.470 177.430 46.695 177.570 ;
        RECT 45.470 177.370 45.790 177.430 ;
        RECT 46.405 177.385 46.695 177.430 ;
        RECT 47.325 177.385 47.615 177.615 ;
        RECT 30.290 177.230 30.610 177.290 ;
        RECT 26.700 177.090 30.610 177.230 ;
        RECT 30.290 177.030 30.610 177.090 ;
        RECT 35.350 177.030 35.670 177.290 ;
        RECT 36.730 177.030 37.050 177.290 ;
        RECT 38.110 177.030 38.430 177.290 ;
        RECT 39.045 177.045 39.335 177.275 ;
        RECT 30.865 176.890 31.155 176.935 ;
        RECT 33.985 176.890 34.275 176.935 ;
        RECT 35.875 176.890 36.165 176.935 ;
        RECT 30.865 176.750 36.165 176.890 ;
        RECT 30.865 176.705 31.155 176.750 ;
        RECT 33.985 176.705 34.275 176.750 ;
        RECT 35.875 176.705 36.165 176.750 ;
        RECT 27.990 176.350 28.310 176.610 ;
        RECT 34.430 176.550 34.750 176.610 ;
        RECT 39.120 176.550 39.260 177.045 ;
        RECT 46.480 176.890 46.620 177.385 ;
        RECT 47.770 177.370 48.090 177.630 ;
        RECT 48.245 177.570 48.535 177.615 ;
        RECT 49.150 177.570 49.470 177.630 ;
        RECT 48.245 177.430 49.470 177.570 ;
        RECT 48.245 177.385 48.535 177.430 ;
        RECT 49.150 177.370 49.470 177.430 ;
        RECT 50.530 177.370 50.850 177.630 ;
        RECT 49.240 177.230 49.380 177.370 ;
        RECT 54.760 177.230 54.900 178.110 ;
        RECT 55.245 177.910 55.535 177.955 ;
        RECT 56.050 177.910 56.370 177.970 ;
        RECT 58.485 177.910 59.135 177.955 ;
        RECT 55.245 177.770 59.135 177.910 ;
        RECT 55.245 177.725 55.835 177.770 ;
        RECT 55.545 177.410 55.835 177.725 ;
        RECT 56.050 177.710 56.370 177.770 ;
        RECT 58.485 177.725 59.135 177.770 ;
        RECT 61.110 177.710 61.430 177.970 ;
        RECT 61.660 177.910 61.800 178.110 ;
        RECT 62.030 178.110 63.715 178.250 ;
        RECT 62.030 178.050 62.350 178.110 ;
        RECT 63.425 178.065 63.715 178.110 ;
        RECT 70.400 178.110 72.455 178.250 ;
        RECT 70.400 177.910 70.540 178.110 ;
        RECT 71.690 178.050 72.010 178.110 ;
        RECT 72.165 178.065 72.455 178.110 ;
        RECT 73.070 178.050 73.390 178.310 ;
        RECT 81.810 178.250 82.130 178.310 ;
        RECT 81.440 178.110 82.130 178.250 ;
        RECT 61.660 177.770 70.540 177.910 ;
        RECT 79.510 177.910 79.830 177.970 ;
        RECT 79.985 177.910 80.275 177.955 ;
        RECT 81.440 177.910 81.580 178.110 ;
        RECT 81.810 178.050 82.130 178.110 ;
        RECT 82.270 178.250 82.590 178.310 ;
        RECT 88.265 178.250 88.555 178.295 ;
        RECT 90.550 178.250 90.870 178.310 ;
        RECT 82.270 178.110 88.020 178.250 ;
        RECT 82.270 178.050 82.590 178.110 ;
        RECT 85.950 177.910 86.270 177.970 ;
        RECT 79.510 177.770 80.275 177.910 ;
        RECT 79.510 177.710 79.830 177.770 ;
        RECT 79.985 177.725 80.275 177.770 ;
        RECT 80.520 177.770 81.580 177.910 ;
        RECT 56.625 177.570 56.915 177.615 ;
        RECT 60.205 177.570 60.495 177.615 ;
        RECT 62.040 177.570 62.330 177.615 ;
        RECT 56.625 177.430 62.330 177.570 ;
        RECT 56.625 177.385 56.915 177.430 ;
        RECT 60.205 177.385 60.495 177.430 ;
        RECT 62.040 177.385 62.330 177.430 ;
        RECT 64.345 177.385 64.635 177.615 ;
        RECT 49.240 177.090 54.900 177.230 ;
        RECT 59.270 177.230 59.590 177.290 ;
        RECT 62.505 177.230 62.795 177.275 ;
        RECT 63.870 177.230 64.190 177.290 ;
        RECT 59.270 177.090 64.190 177.230 ;
        RECT 59.270 177.030 59.590 177.090 ;
        RECT 62.505 177.045 62.795 177.090 ;
        RECT 63.870 177.030 64.190 177.090 ;
        RECT 50.990 176.890 51.310 176.950 ;
        RECT 46.480 176.750 51.310 176.890 ;
        RECT 50.990 176.690 51.310 176.750 ;
        RECT 56.625 176.890 56.915 176.935 ;
        RECT 59.745 176.890 60.035 176.935 ;
        RECT 61.635 176.890 61.925 176.935 ;
        RECT 56.625 176.750 61.925 176.890 ;
        RECT 56.625 176.705 56.915 176.750 ;
        RECT 59.745 176.705 60.035 176.750 ;
        RECT 61.635 176.705 61.925 176.750 ;
        RECT 34.430 176.410 39.260 176.550 ;
        RECT 41.345 176.550 41.635 176.595 ;
        RECT 42.710 176.550 43.030 176.610 ;
        RECT 41.345 176.410 43.030 176.550 ;
        RECT 34.430 176.350 34.750 176.410 ;
        RECT 41.345 176.365 41.635 176.410 ;
        RECT 42.710 176.350 43.030 176.410 ;
        RECT 49.625 176.550 49.915 176.595 ;
        RECT 50.070 176.550 50.390 176.610 ;
        RECT 49.625 176.410 50.390 176.550 ;
        RECT 49.625 176.365 49.915 176.410 ;
        RECT 50.070 176.350 50.390 176.410 ;
        RECT 53.305 176.550 53.595 176.595 ;
        RECT 64.420 176.550 64.560 177.385 ;
        RECT 68.930 177.370 69.250 177.630 ;
        RECT 69.390 177.570 69.710 177.630 ;
        RECT 71.280 177.570 71.570 177.615 ;
        RECT 72.610 177.570 72.930 177.630 ;
        RECT 73.545 177.570 73.835 177.615 ;
        RECT 69.390 177.430 72.380 177.570 ;
        RECT 69.390 177.370 69.710 177.430 ;
        RECT 71.280 177.385 71.570 177.430 ;
        RECT 72.240 177.230 72.380 177.430 ;
        RECT 72.610 177.430 73.835 177.570 ;
        RECT 72.610 177.370 72.930 177.430 ;
        RECT 73.545 177.385 73.835 177.430 ;
        RECT 73.990 177.370 74.310 177.630 ;
        RECT 74.910 177.370 75.230 177.630 ;
        RECT 75.385 177.385 75.675 177.615 ;
        RECT 75.460 177.230 75.600 177.385 ;
        RECT 76.290 177.370 76.610 177.630 ;
        RECT 77.225 177.385 77.515 177.615 ;
        RECT 72.240 177.090 75.600 177.230 ;
        RECT 77.300 177.230 77.440 177.385 ;
        RECT 77.670 177.370 77.990 177.630 ;
        RECT 78.130 177.570 78.450 177.630 ;
        RECT 80.520 177.570 80.660 177.770 ;
        RECT 81.440 177.615 81.580 177.770 ;
        RECT 82.360 177.770 86.270 177.910 ;
        RECT 87.880 177.910 88.020 178.110 ;
        RECT 88.265 178.110 90.870 178.250 ;
        RECT 88.265 178.065 88.555 178.110 ;
        RECT 90.550 178.050 90.870 178.110 ;
        RECT 99.750 178.250 100.070 178.310 ;
        RECT 102.065 178.250 102.355 178.295 ;
        RECT 99.750 178.110 102.355 178.250 ;
        RECT 99.750 178.050 100.070 178.110 ;
        RECT 102.065 178.065 102.355 178.110 ;
        RECT 111.710 178.050 112.030 178.310 ;
        RECT 112.170 178.050 112.490 178.310 ;
        RECT 114.025 178.065 114.315 178.295 ;
        RECT 117.705 178.250 117.995 178.295 ;
        RECT 118.610 178.250 118.930 178.310 ;
        RECT 117.705 178.110 118.930 178.250 ;
        RECT 117.705 178.065 117.995 178.110 ;
        RECT 108.950 177.910 109.270 177.970 ;
        RECT 87.880 177.770 106.880 177.910 ;
        RECT 78.130 177.430 80.660 177.570 ;
        RECT 78.130 177.370 78.450 177.430 ;
        RECT 81.365 177.385 81.655 177.615 ;
        RECT 81.810 177.370 82.130 177.630 ;
        RECT 82.360 177.615 82.500 177.770 ;
        RECT 85.950 177.710 86.270 177.770 ;
        RECT 82.285 177.385 82.575 177.615 ;
        RECT 82.730 177.570 83.050 177.630 ;
        RECT 83.205 177.570 83.495 177.615 ;
        RECT 84.110 177.570 84.430 177.630 ;
        RECT 82.730 177.430 84.430 177.570 ;
        RECT 82.730 177.370 83.050 177.430 ;
        RECT 83.205 177.385 83.495 177.430 ;
        RECT 84.110 177.370 84.430 177.430 ;
        RECT 85.505 177.570 85.795 177.615 ;
        RECT 89.170 177.570 89.490 177.630 ;
        RECT 85.505 177.430 89.490 177.570 ;
        RECT 85.505 177.385 85.795 177.430 ;
        RECT 89.170 177.370 89.490 177.430 ;
        RECT 98.370 177.370 98.690 177.630 ;
        RECT 99.290 177.370 99.610 177.630 ;
        RECT 99.840 177.615 99.980 177.770 ;
        RECT 106.740 177.630 106.880 177.770 ;
        RECT 107.200 177.770 109.270 177.910 ;
        RECT 114.100 177.910 114.240 178.065 ;
        RECT 118.610 178.050 118.930 178.110 ;
        RECT 121.830 177.910 122.150 177.970 ;
        RECT 114.100 177.770 122.150 177.910 ;
        RECT 99.765 177.385 100.055 177.615 ;
        RECT 100.225 177.385 100.515 177.615 ;
        RECT 102.050 177.570 102.370 177.630 ;
        RECT 102.985 177.570 103.275 177.615 ;
        RECT 102.050 177.430 103.275 177.570 ;
        RECT 79.050 177.230 79.370 177.290 ;
        RECT 77.300 177.090 79.370 177.230 ;
        RECT 79.050 177.030 79.370 177.090 ;
        RECT 79.525 177.230 79.815 177.275 ;
        RECT 80.430 177.230 80.750 177.290 ;
        RECT 100.300 177.230 100.440 177.385 ;
        RECT 102.050 177.370 102.370 177.430 ;
        RECT 102.985 177.385 103.275 177.430 ;
        RECT 106.205 177.385 106.495 177.615 ;
        RECT 105.730 177.230 106.050 177.290 ;
        RECT 106.280 177.230 106.420 177.385 ;
        RECT 106.650 177.370 106.970 177.630 ;
        RECT 107.200 177.615 107.340 177.770 ;
        RECT 108.950 177.710 109.270 177.770 ;
        RECT 121.830 177.710 122.150 177.770 ;
        RECT 107.125 177.385 107.415 177.615 ;
        RECT 108.030 177.570 108.350 177.630 ;
        RECT 109.410 177.570 109.730 177.630 ;
        RECT 108.030 177.430 109.730 177.570 ;
        RECT 108.030 177.370 108.350 177.430 ;
        RECT 109.410 177.370 109.730 177.430 ;
        RECT 116.770 177.370 117.090 177.630 ;
        RECT 79.525 177.090 80.750 177.230 ;
        RECT 79.525 177.045 79.815 177.090 ;
        RECT 80.430 177.030 80.750 177.090 ;
        RECT 84.890 177.090 106.420 177.230 ;
        RECT 65.250 176.890 65.570 176.950 ;
        RECT 70.325 176.890 70.615 176.935 ;
        RECT 84.890 176.890 85.030 177.090 ;
        RECT 105.730 177.030 106.050 177.090 ;
        RECT 110.790 177.030 111.110 177.290 ;
        RECT 65.250 176.750 85.030 176.890 ;
        RECT 65.250 176.690 65.570 176.750 ;
        RECT 70.325 176.705 70.615 176.750 ;
        RECT 53.305 176.410 64.560 176.550 ;
        RECT 64.790 176.550 65.110 176.610 ;
        RECT 68.010 176.550 68.330 176.610 ;
        RECT 64.790 176.410 68.330 176.550 ;
        RECT 53.305 176.365 53.595 176.410 ;
        RECT 64.790 176.350 65.110 176.410 ;
        RECT 68.010 176.350 68.330 176.410 ;
        RECT 68.930 176.550 69.250 176.610 ;
        RECT 74.910 176.550 75.230 176.610 ;
        RECT 68.930 176.410 75.230 176.550 ;
        RECT 68.930 176.350 69.250 176.410 ;
        RECT 74.910 176.350 75.230 176.410 ;
        RECT 100.670 176.550 100.990 176.610 ;
        RECT 101.605 176.550 101.895 176.595 ;
        RECT 100.670 176.410 101.895 176.550 ;
        RECT 100.670 176.350 100.990 176.410 ;
        RECT 101.605 176.365 101.895 176.410 ;
        RECT 102.050 176.550 102.370 176.610 ;
        RECT 104.825 176.550 105.115 176.595 ;
        RECT 102.050 176.410 105.115 176.550 ;
        RECT 102.050 176.350 102.370 176.410 ;
        RECT 104.825 176.365 105.115 176.410 ;
        RECT 14.580 175.730 127.740 176.210 ;
        RECT 25.705 175.530 25.995 175.575 ;
        RECT 26.150 175.530 26.470 175.590 ;
        RECT 38.110 175.530 38.430 175.590 ;
        RECT 40.870 175.530 41.190 175.590 ;
        RECT 25.705 175.390 26.470 175.530 ;
        RECT 25.705 175.345 25.995 175.390 ;
        RECT 26.150 175.330 26.470 175.390 ;
        RECT 34.060 175.390 38.430 175.530 ;
        RECT 30.765 175.190 31.055 175.235 ;
        RECT 26.700 175.050 31.055 175.190 ;
        RECT 26.700 174.555 26.840 175.050 ;
        RECT 30.765 175.005 31.055 175.050 ;
        RECT 34.060 174.895 34.200 175.390 ;
        RECT 38.110 175.330 38.430 175.390 ;
        RECT 38.660 175.390 41.190 175.530 ;
        RECT 38.660 175.190 38.800 175.390 ;
        RECT 40.870 175.330 41.190 175.390 ;
        RECT 46.390 175.530 46.710 175.590 ;
        RECT 54.210 175.530 54.530 175.590 ;
        RECT 46.390 175.390 54.530 175.530 ;
        RECT 46.390 175.330 46.710 175.390 ;
        RECT 54.210 175.330 54.530 175.390 ;
        RECT 63.870 175.530 64.190 175.590 ;
        RECT 66.170 175.530 66.490 175.590 ;
        RECT 63.870 175.390 66.490 175.530 ;
        RECT 63.870 175.330 64.190 175.390 ;
        RECT 66.170 175.330 66.490 175.390 ;
        RECT 68.010 175.530 68.330 175.590 ;
        RECT 77.670 175.530 77.990 175.590 ;
        RECT 81.810 175.530 82.130 175.590 ;
        RECT 106.190 175.530 106.510 175.590 ;
        RECT 108.030 175.530 108.350 175.590 ;
        RECT 68.010 175.390 82.130 175.530 ;
        RECT 68.010 175.330 68.330 175.390 ;
        RECT 77.670 175.330 77.990 175.390 ;
        RECT 81.810 175.330 82.130 175.390 ;
        RECT 103.980 175.390 110.560 175.530 ;
        RECT 36.820 175.050 38.800 175.190 ;
        RECT 39.045 175.190 39.335 175.235 ;
        RECT 40.410 175.190 40.730 175.250 ;
        RECT 57.445 175.190 57.735 175.235 ;
        RECT 39.045 175.050 40.730 175.190 ;
        RECT 33.985 174.665 34.275 174.895 ;
        RECT 36.820 174.850 36.960 175.050 ;
        RECT 39.045 175.005 39.335 175.050 ;
        RECT 40.410 174.990 40.730 175.050 ;
        RECT 53.840 175.050 57.735 175.190 ;
        RECT 53.840 174.910 53.980 175.050 ;
        RECT 57.445 175.005 57.735 175.050 ;
        RECT 60.305 175.190 60.595 175.235 ;
        RECT 63.425 175.190 63.715 175.235 ;
        RECT 65.315 175.190 65.605 175.235 ;
        RECT 71.705 175.190 71.995 175.235 ;
        RECT 76.290 175.190 76.610 175.250 ;
        RECT 60.305 175.050 65.605 175.190 ;
        RECT 60.305 175.005 60.595 175.050 ;
        RECT 63.425 175.005 63.715 175.050 ;
        RECT 65.315 175.005 65.605 175.050 ;
        RECT 69.480 175.050 76.610 175.190 ;
        RECT 35.440 174.710 36.960 174.850 ;
        RECT 37.650 174.850 37.970 174.910 ;
        RECT 45.470 174.850 45.790 174.910 ;
        RECT 37.650 174.710 41.560 174.850 ;
        RECT 26.625 174.325 26.915 174.555 ;
        RECT 27.085 174.325 27.375 174.555 ;
        RECT 30.305 174.510 30.595 174.555 ;
        RECT 32.605 174.510 32.895 174.555 ;
        RECT 34.430 174.510 34.750 174.570 ;
        RECT 35.440 174.555 35.580 174.710 ;
        RECT 37.650 174.650 37.970 174.710 ;
        RECT 30.305 174.370 34.750 174.510 ;
        RECT 30.305 174.325 30.595 174.370 ;
        RECT 32.605 174.325 32.895 174.370 ;
        RECT 27.160 174.170 27.300 174.325 ;
        RECT 34.430 174.310 34.750 174.370 ;
        RECT 35.365 174.325 35.655 174.555 ;
        RECT 36.285 174.325 36.575 174.555 ;
        RECT 36.745 174.325 37.035 174.555 ;
        RECT 37.205 174.510 37.495 174.555 ;
        RECT 38.110 174.510 38.430 174.570 ;
        RECT 39.950 174.510 40.270 174.570 ;
        RECT 41.420 174.555 41.560 174.710 ;
        RECT 42.800 174.710 45.790 174.850 ;
        RECT 42.800 174.555 42.940 174.710 ;
        RECT 45.470 174.650 45.790 174.710 ;
        RECT 46.865 174.850 47.155 174.895 ;
        RECT 53.750 174.850 54.070 174.910 ;
        RECT 46.865 174.710 54.070 174.850 ;
        RECT 46.865 174.665 47.155 174.710 ;
        RECT 53.750 174.650 54.070 174.710 ;
        RECT 54.210 174.650 54.530 174.910 ;
        RECT 57.890 174.850 58.210 174.910 ;
        RECT 64.790 174.850 65.110 174.910 ;
        RECT 54.760 174.710 58.210 174.850 ;
        RECT 40.425 174.510 40.715 174.555 ;
        RECT 37.205 174.370 40.715 174.510 ;
        RECT 37.205 174.325 37.495 174.370 ;
        RECT 27.990 174.170 28.310 174.230 ;
        RECT 33.065 174.170 33.355 174.215 ;
        RECT 33.970 174.170 34.290 174.230 ;
        RECT 36.360 174.170 36.500 174.325 ;
        RECT 27.160 174.030 32.820 174.170 ;
        RECT 27.990 173.970 28.310 174.030 ;
        RECT 32.680 173.830 32.820 174.030 ;
        RECT 33.065 174.030 34.290 174.170 ;
        RECT 33.065 173.985 33.355 174.030 ;
        RECT 33.970 173.970 34.290 174.030 ;
        RECT 34.520 174.030 36.500 174.170 ;
        RECT 34.520 173.830 34.660 174.030 ;
        RECT 32.680 173.690 34.660 173.830 ;
        RECT 36.820 173.830 36.960 174.325 ;
        RECT 38.110 174.310 38.430 174.370 ;
        RECT 39.950 174.310 40.270 174.370 ;
        RECT 40.425 174.325 40.715 174.370 ;
        RECT 40.885 174.325 41.175 174.555 ;
        RECT 41.345 174.325 41.635 174.555 ;
        RECT 42.265 174.510 42.555 174.555 ;
        RECT 42.725 174.510 43.015 174.555 ;
        RECT 42.265 174.370 43.015 174.510 ;
        RECT 42.265 174.325 42.555 174.370 ;
        RECT 42.725 174.325 43.015 174.370 ;
        RECT 38.585 174.170 38.875 174.215 ;
        RECT 39.030 174.170 39.350 174.230 ;
        RECT 38.585 174.030 39.350 174.170 ;
        RECT 38.585 173.985 38.875 174.030 ;
        RECT 39.030 173.970 39.350 174.030 ;
        RECT 39.490 174.170 39.810 174.230 ;
        RECT 40.960 174.170 41.100 174.325 ;
        RECT 43.630 174.310 43.950 174.570 ;
        RECT 44.090 174.310 44.410 174.570 ;
        RECT 44.550 174.310 44.870 174.570 ;
        RECT 54.760 174.555 54.900 174.710 ;
        RECT 57.890 174.650 58.210 174.710 ;
        RECT 58.440 174.710 65.110 174.850 ;
        RECT 49.625 174.510 49.915 174.555 ;
        RECT 54.685 174.510 54.975 174.555 ;
        RECT 49.625 174.370 54.975 174.510 ;
        RECT 49.625 174.325 49.915 174.370 ;
        RECT 54.685 174.325 54.975 174.370 ;
        RECT 55.145 174.510 55.435 174.555 ;
        RECT 56.510 174.510 56.830 174.570 ;
        RECT 55.145 174.370 56.830 174.510 ;
        RECT 55.145 174.325 55.435 174.370 ;
        RECT 56.510 174.310 56.830 174.370 ;
        RECT 41.790 174.170 42.110 174.230 ;
        RECT 39.490 174.030 42.110 174.170 ;
        RECT 39.490 173.970 39.810 174.030 ;
        RECT 41.790 173.970 42.110 174.030 ;
        RECT 39.580 173.830 39.720 173.970 ;
        RECT 36.820 173.690 39.720 173.830 ;
        RECT 44.180 173.830 44.320 174.310 ;
        RECT 45.470 174.170 45.790 174.230 ;
        RECT 45.945 174.170 46.235 174.215 ;
        RECT 45.470 174.030 46.235 174.170 ;
        RECT 45.470 173.970 45.790 174.030 ;
        RECT 45.945 173.985 46.235 174.030 ;
        RECT 47.770 174.170 48.090 174.230 ;
        RECT 53.290 174.170 53.610 174.230 ;
        RECT 58.440 174.170 58.580 174.710 ;
        RECT 64.790 174.650 65.110 174.710 ;
        RECT 66.170 174.650 66.490 174.910 ;
        RECT 59.225 174.215 59.515 174.530 ;
        RECT 60.305 174.510 60.595 174.555 ;
        RECT 63.885 174.510 64.175 174.555 ;
        RECT 65.720 174.510 66.010 174.555 ;
        RECT 60.305 174.370 66.010 174.510 ;
        RECT 60.305 174.325 60.595 174.370 ;
        RECT 63.885 174.325 64.175 174.370 ;
        RECT 65.720 174.325 66.010 174.370 ;
        RECT 68.485 174.510 68.775 174.555 ;
        RECT 68.930 174.510 69.250 174.570 ;
        RECT 68.485 174.370 69.250 174.510 ;
        RECT 68.485 174.325 68.775 174.370 ;
        RECT 68.930 174.310 69.250 174.370 ;
        RECT 47.770 174.030 58.580 174.170 ;
        RECT 58.925 174.170 59.515 174.215 ;
        RECT 61.110 174.170 61.430 174.230 ;
        RECT 62.165 174.170 62.815 174.215 ;
        RECT 58.925 174.030 62.815 174.170 ;
        RECT 47.770 173.970 48.090 174.030 ;
        RECT 53.290 173.970 53.610 174.030 ;
        RECT 58.925 173.985 59.215 174.030 ;
        RECT 61.110 173.970 61.430 174.030 ;
        RECT 62.165 173.985 62.815 174.030 ;
        RECT 64.790 173.970 65.110 174.230 ;
        RECT 69.480 174.170 69.620 175.050 ;
        RECT 71.705 175.005 71.995 175.050 ;
        RECT 76.290 174.990 76.610 175.050 ;
        RECT 69.850 174.650 70.170 174.910 ;
        RECT 81.900 174.850 82.040 175.330 ;
        RECT 87.330 174.850 87.650 174.910 ;
        RECT 81.900 174.710 82.960 174.850 ;
        RECT 72.610 174.310 72.930 174.570 ;
        RECT 78.130 174.510 78.450 174.570 ;
        RECT 82.820 174.555 82.960 174.710 ;
        RECT 83.280 174.710 87.650 174.850 ;
        RECT 83.280 174.555 83.420 174.710 ;
        RECT 87.330 174.650 87.650 174.710 ;
        RECT 82.285 174.510 82.575 174.555 ;
        RECT 78.130 174.370 82.575 174.510 ;
        RECT 78.130 174.310 78.450 174.370 ;
        RECT 82.285 174.325 82.575 174.370 ;
        RECT 82.745 174.325 83.035 174.555 ;
        RECT 83.205 174.325 83.495 174.555 ;
        RECT 84.110 174.310 84.430 174.570 ;
        RECT 98.370 174.510 98.690 174.570 ;
        RECT 103.980 174.555 104.120 175.390 ;
        RECT 106.190 175.330 106.510 175.390 ;
        RECT 108.030 175.330 108.350 175.390 ;
        RECT 107.125 175.190 107.415 175.235 ;
        RECT 108.950 175.190 109.270 175.250 ;
        RECT 107.125 175.050 109.270 175.190 ;
        RECT 107.125 175.005 107.415 175.050 ;
        RECT 108.950 174.990 109.270 175.050 ;
        RECT 106.650 174.850 106.970 174.910 ;
        RECT 105.360 174.710 109.640 174.850 ;
        RECT 103.905 174.510 104.195 174.555 ;
        RECT 98.370 174.370 104.195 174.510 ;
        RECT 98.370 174.310 98.690 174.370 ;
        RECT 103.905 174.325 104.195 174.370 ;
        RECT 104.810 174.310 105.130 174.570 ;
        RECT 105.360 174.555 105.500 174.710 ;
        RECT 106.650 174.650 106.970 174.710 ;
        RECT 109.500 174.570 109.640 174.710 ;
        RECT 105.285 174.325 105.575 174.555 ;
        RECT 105.730 174.510 106.050 174.570 ;
        RECT 108.965 174.510 109.255 174.555 ;
        RECT 105.730 174.370 109.255 174.510 ;
        RECT 105.730 174.310 106.050 174.370 ;
        RECT 108.965 174.325 109.255 174.370 ;
        RECT 65.340 174.030 69.620 174.170 ;
        RECT 80.905 174.170 81.195 174.215 ;
        RECT 81.810 174.170 82.130 174.230 ;
        RECT 80.905 174.030 82.130 174.170 ;
        RECT 47.860 173.830 48.000 173.970 ;
        RECT 44.180 173.690 48.000 173.830 ;
        RECT 56.970 173.630 57.290 173.890 ;
        RECT 62.950 173.830 63.270 173.890 ;
        RECT 65.340 173.830 65.480 174.030 ;
        RECT 80.905 173.985 81.195 174.030 ;
        RECT 81.810 173.970 82.130 174.030 ;
        RECT 104.350 174.170 104.670 174.230 ;
        RECT 107.585 174.170 107.875 174.215 ;
        RECT 104.350 174.030 107.875 174.170 ;
        RECT 104.350 173.970 104.670 174.030 ;
        RECT 107.585 173.985 107.875 174.030 ;
        RECT 62.950 173.690 65.480 173.830 ;
        RECT 70.770 173.830 71.090 173.890 ;
        RECT 98.370 173.830 98.690 173.890 ;
        RECT 70.770 173.690 98.690 173.830 ;
        RECT 109.040 173.830 109.180 174.325 ;
        RECT 109.410 174.310 109.730 174.570 ;
        RECT 109.870 174.310 110.190 174.570 ;
        RECT 110.420 174.510 110.560 175.390 ;
        RECT 110.805 174.510 111.095 174.555 ;
        RECT 110.420 174.370 111.095 174.510 ;
        RECT 110.805 174.325 111.095 174.370 ;
        RECT 118.165 174.510 118.455 174.555 ;
        RECT 119.070 174.510 119.390 174.570 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 118.165 174.370 119.390 174.510 ;
        RECT 118.165 174.325 118.455 174.370 ;
        RECT 119.070 174.310 119.390 174.370 ;
        RECT 118.625 173.985 118.915 174.215 ;
        RECT 109.870 173.830 110.190 173.890 ;
        RECT 109.040 173.690 110.190 173.830 ;
        RECT 62.950 173.630 63.270 173.690 ;
        RECT 70.770 173.630 71.090 173.690 ;
        RECT 98.370 173.630 98.690 173.690 ;
        RECT 109.870 173.630 110.190 173.690 ;
        RECT 118.150 173.830 118.470 173.890 ;
        RECT 118.700 173.830 118.840 173.985 ;
        RECT 118.150 173.690 118.840 173.830 ;
        RECT 118.150 173.630 118.470 173.690 ;
        RECT 14.580 173.010 127.740 173.490 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 35.350 172.810 35.670 172.870 ;
        RECT 41.805 172.810 42.095 172.855 ;
        RECT 35.350 172.670 42.095 172.810 ;
        RECT 35.350 172.610 35.670 172.670 ;
        RECT 41.805 172.625 42.095 172.670 ;
        RECT 44.550 172.810 44.870 172.870 ;
        RECT 49.150 172.810 49.470 172.870 ;
        RECT 44.550 172.670 49.470 172.810 ;
        RECT 44.550 172.610 44.870 172.670 ;
        RECT 37.190 172.470 37.510 172.530 ;
        RECT 37.190 172.330 40.180 172.470 ;
        RECT 37.190 172.270 37.510 172.330 ;
        RECT 38.110 172.130 38.430 172.190 ;
        RECT 39.045 172.130 39.335 172.175 ;
        RECT 38.110 171.990 39.335 172.130 ;
        RECT 38.110 171.930 38.430 171.990 ;
        RECT 39.045 171.945 39.335 171.990 ;
        RECT 39.490 171.930 39.810 172.190 ;
        RECT 40.040 172.175 40.180 172.330 ;
        RECT 39.965 171.945 40.255 172.175 ;
        RECT 40.870 171.930 41.190 172.190 ;
        RECT 42.710 171.930 43.030 172.190 ;
        RECT 45.560 172.175 45.700 172.670 ;
        RECT 49.150 172.610 49.470 172.670 ;
        RECT 49.610 172.810 49.930 172.870 ;
        RECT 50.990 172.810 51.310 172.870 ;
        RECT 54.670 172.810 54.990 172.870 ;
        RECT 49.610 172.670 50.300 172.810 ;
        RECT 49.610 172.610 49.930 172.670 ;
        RECT 46.020 172.330 49.840 172.470 ;
        RECT 46.020 172.175 46.160 172.330 ;
        RECT 49.700 172.190 49.840 172.330 ;
        RECT 45.485 171.945 45.775 172.175 ;
        RECT 45.945 171.945 46.235 172.175 ;
        RECT 46.405 171.945 46.695 172.175 ;
        RECT 35.810 171.790 36.130 171.850 ;
        RECT 46.480 171.790 46.620 171.945 ;
        RECT 47.310 171.930 47.630 172.190 ;
        RECT 49.150 171.930 49.470 172.190 ;
        RECT 49.610 171.930 49.930 172.190 ;
        RECT 50.160 172.175 50.300 172.670 ;
        RECT 50.990 172.670 54.990 172.810 ;
        RECT 50.990 172.610 51.310 172.670 ;
        RECT 54.670 172.610 54.990 172.670 ;
        RECT 60.665 172.810 60.955 172.855 ;
        RECT 61.110 172.810 61.430 172.870 ;
        RECT 60.665 172.670 61.430 172.810 ;
        RECT 60.665 172.625 60.955 172.670 ;
        RECT 61.110 172.610 61.430 172.670 ;
        RECT 62.505 172.810 62.795 172.855 ;
        RECT 64.790 172.810 65.110 172.870 ;
        RECT 91.010 172.810 91.330 172.870 ;
        RECT 119.070 172.810 119.390 172.870 ;
        RECT 62.505 172.670 65.110 172.810 ;
        RECT 62.505 172.625 62.795 172.670 ;
        RECT 64.790 172.610 65.110 172.670 ;
        RECT 89.720 172.670 99.980 172.810 ;
        RECT 56.970 172.470 57.290 172.530 ;
        RECT 83.665 172.470 83.955 172.515 ;
        RECT 89.720 172.470 89.860 172.670 ;
        RECT 91.010 172.610 91.330 172.670 ;
        RECT 56.970 172.330 61.800 172.470 ;
        RECT 56.970 172.270 57.290 172.330 ;
        RECT 50.085 171.945 50.375 172.175 ;
        RECT 50.990 171.930 51.310 172.190 ;
        RECT 52.845 171.945 53.135 172.175 ;
        RECT 35.810 171.650 46.620 171.790 ;
        RECT 49.240 171.790 49.380 171.930 ;
        RECT 52.920 171.790 53.060 171.945 ;
        RECT 53.290 171.930 53.610 172.190 ;
        RECT 53.750 171.930 54.070 172.190 ;
        RECT 54.670 171.930 54.990 172.190 ;
        RECT 60.650 172.130 60.970 172.190 ;
        RECT 61.660 172.175 61.800 172.330 ;
        RECT 83.665 172.330 89.860 172.470 ;
        RECT 83.665 172.285 83.955 172.330 ;
        RECT 61.125 172.130 61.415 172.175 ;
        RECT 60.650 171.990 61.415 172.130 ;
        RECT 60.650 171.930 60.970 171.990 ;
        RECT 61.125 171.945 61.415 171.990 ;
        RECT 61.585 171.945 61.875 172.175 ;
        RECT 68.930 172.130 69.250 172.190 ;
        RECT 89.720 172.175 89.860 172.330 ;
        RECT 90.105 172.470 90.395 172.515 ;
        RECT 92.505 172.470 92.795 172.515 ;
        RECT 95.745 172.470 96.395 172.515 ;
        RECT 90.105 172.330 96.395 172.470 ;
        RECT 90.105 172.285 90.395 172.330 ;
        RECT 92.505 172.285 93.095 172.330 ;
        RECT 95.745 172.285 96.395 172.330 ;
        RECT 82.285 172.130 82.575 172.175 ;
        RECT 68.930 171.990 82.575 172.130 ;
        RECT 68.930 171.930 69.250 171.990 ;
        RECT 82.285 171.945 82.575 171.990 ;
        RECT 89.645 171.945 89.935 172.175 ;
        RECT 92.805 171.970 93.095 172.285 ;
        RECT 93.885 172.130 94.175 172.175 ;
        RECT 97.465 172.130 97.755 172.175 ;
        RECT 99.300 172.130 99.590 172.175 ;
        RECT 93.885 171.990 99.590 172.130 ;
        RECT 99.840 172.130 99.980 172.670 ;
        RECT 113.180 172.670 119.390 172.810 ;
        RECT 106.190 172.470 106.510 172.530 ;
        RECT 110.330 172.470 110.650 172.530 ;
        RECT 106.190 172.330 108.260 172.470 ;
        RECT 106.190 172.270 106.510 172.330 ;
        RECT 108.120 172.175 108.260 172.330 ;
        RECT 109.040 172.330 110.650 172.470 ;
        RECT 109.040 172.175 109.180 172.330 ;
        RECT 110.330 172.270 110.650 172.330 ;
        RECT 107.585 172.130 107.875 172.175 ;
        RECT 99.840 171.990 107.875 172.130 ;
        RECT 93.885 171.945 94.175 171.990 ;
        RECT 97.465 171.945 97.755 171.990 ;
        RECT 99.300 171.945 99.590 171.990 ;
        RECT 107.585 171.945 107.875 171.990 ;
        RECT 108.045 171.945 108.335 172.175 ;
        RECT 108.965 171.945 109.255 172.175 ;
        RECT 49.240 171.650 53.060 171.790 ;
        RECT 35.810 171.590 36.130 171.650 ;
        RECT 49.610 171.450 49.930 171.510 ;
        RECT 53.380 171.450 53.520 171.930 ;
        RECT 85.505 171.790 85.795 171.835 ;
        RECT 85.505 171.650 91.240 171.790 ;
        RECT 85.505 171.605 85.795 171.650 ;
        RECT 49.610 171.310 53.520 171.450 ;
        RECT 49.610 171.250 49.930 171.310 ;
        RECT 35.350 171.110 35.670 171.170 ;
        RECT 37.665 171.110 37.955 171.155 ;
        RECT 35.350 170.970 37.955 171.110 ;
        RECT 35.350 170.910 35.670 170.970 ;
        RECT 37.665 170.925 37.955 170.970 ;
        RECT 41.330 171.110 41.650 171.170 ;
        RECT 44.105 171.110 44.395 171.155 ;
        RECT 41.330 170.970 44.395 171.110 ;
        RECT 41.330 170.910 41.650 170.970 ;
        RECT 44.105 170.925 44.395 170.970 ;
        RECT 45.930 171.110 46.250 171.170 ;
        RECT 47.785 171.110 48.075 171.155 ;
        RECT 45.930 170.970 48.075 171.110 ;
        RECT 45.930 170.910 46.250 170.970 ;
        RECT 47.785 170.925 48.075 170.970 ;
        RECT 51.465 171.110 51.755 171.155 ;
        RECT 52.370 171.110 52.690 171.170 ;
        RECT 51.465 170.970 52.690 171.110 ;
        RECT 51.465 170.925 51.755 170.970 ;
        RECT 52.370 170.910 52.690 170.970 ;
        RECT 88.265 171.110 88.555 171.155 ;
        RECT 89.630 171.110 89.950 171.170 ;
        RECT 91.100 171.155 91.240 171.650 ;
        RECT 98.370 171.590 98.690 171.850 ;
        RECT 99.765 171.790 100.055 171.835 ;
        RECT 105.730 171.790 106.050 171.850 ;
        RECT 99.765 171.650 106.050 171.790 ;
        RECT 107.660 171.790 107.800 171.945 ;
        RECT 109.410 171.930 109.730 172.190 ;
        RECT 109.870 171.930 110.190 172.190 ;
        RECT 113.180 172.175 113.320 172.670 ;
        RECT 119.070 172.610 119.390 172.670 ;
        RECT 117.345 172.470 117.635 172.515 ;
        RECT 118.150 172.470 118.470 172.530 ;
        RECT 120.585 172.470 121.235 172.515 ;
        RECT 117.345 172.330 121.235 172.470 ;
        RECT 117.345 172.285 117.935 172.330 ;
        RECT 113.105 171.945 113.395 172.175 ;
        RECT 117.645 171.970 117.935 172.285 ;
        RECT 118.150 172.270 118.470 172.330 ;
        RECT 120.585 172.285 121.235 172.330 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 118.725 172.130 119.015 172.175 ;
        RECT 122.305 172.130 122.595 172.175 ;
        RECT 124.140 172.130 124.430 172.175 ;
        RECT 118.725 171.990 124.430 172.130 ;
        RECT 118.725 171.945 119.015 171.990 ;
        RECT 122.305 171.945 122.595 171.990 ;
        RECT 124.140 171.945 124.430 171.990 ;
        RECT 113.180 171.790 113.320 171.945 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 107.660 171.650 113.320 171.790 ;
        RECT 121.370 171.790 121.690 171.850 ;
        RECT 123.225 171.790 123.515 171.835 ;
        RECT 121.370 171.650 123.515 171.790 ;
        RECT 99.765 171.605 100.055 171.650 ;
        RECT 105.730 171.590 106.050 171.650 ;
        RECT 121.370 171.590 121.690 171.650 ;
        RECT 123.225 171.605 123.515 171.650 ;
        RECT 124.590 171.590 124.910 171.850 ;
        RECT 93.885 171.450 94.175 171.495 ;
        RECT 97.005 171.450 97.295 171.495 ;
        RECT 98.895 171.450 99.185 171.495 ;
        RECT 114.470 171.450 114.790 171.510 ;
        RECT 93.885 171.310 99.185 171.450 ;
        RECT 93.885 171.265 94.175 171.310 ;
        RECT 97.005 171.265 97.295 171.310 ;
        RECT 98.895 171.265 99.185 171.310 ;
        RECT 99.840 171.310 114.790 171.450 ;
        RECT 88.265 170.970 89.950 171.110 ;
        RECT 88.265 170.925 88.555 170.970 ;
        RECT 89.630 170.910 89.950 170.970 ;
        RECT 91.025 171.110 91.315 171.155 ;
        RECT 99.840 171.110 99.980 171.310 ;
        RECT 114.470 171.250 114.790 171.310 ;
        RECT 118.725 171.450 119.015 171.495 ;
        RECT 121.845 171.450 122.135 171.495 ;
        RECT 123.735 171.450 124.025 171.495 ;
        RECT 118.725 171.310 124.025 171.450 ;
        RECT 118.725 171.265 119.015 171.310 ;
        RECT 121.845 171.265 122.135 171.310 ;
        RECT 123.735 171.265 124.025 171.310 ;
        RECT 91.025 170.970 99.980 171.110 ;
        RECT 91.025 170.925 91.315 170.970 ;
        RECT 107.110 170.910 107.430 171.170 ;
        RECT 111.250 170.910 111.570 171.170 ;
        RECT 113.550 170.910 113.870 171.170 ;
        RECT 115.865 171.110 116.155 171.155 ;
        RECT 117.230 171.110 117.550 171.170 ;
        RECT 115.865 170.970 117.550 171.110 ;
        RECT 115.865 170.925 116.155 170.970 ;
        RECT 117.230 170.910 117.550 170.970 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 14.580 170.290 127.740 170.770 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 47.310 170.090 47.630 170.150 ;
        RECT 67.550 170.090 67.870 170.150 ;
        RECT 68.945 170.090 69.235 170.135 ;
        RECT 47.310 169.950 69.235 170.090 ;
        RECT 47.310 169.890 47.630 169.950 ;
        RECT 67.550 169.890 67.870 169.950 ;
        RECT 68.945 169.905 69.235 169.950 ;
        RECT 70.770 169.890 71.090 170.150 ;
        RECT 97.005 170.090 97.295 170.135 ;
        RECT 98.370 170.090 98.690 170.150 ;
        RECT 97.005 169.950 98.690 170.090 ;
        RECT 97.005 169.905 97.295 169.950 ;
        RECT 98.370 169.890 98.690 169.950 ;
        RECT 121.370 169.890 121.690 170.150 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 40.870 169.750 41.190 169.810 ;
        RECT 70.860 169.750 71.000 169.890 ;
        RECT 40.870 169.610 71.000 169.750 ;
        RECT 84.540 169.750 84.830 169.795 ;
        RECT 87.320 169.750 87.610 169.795 ;
        RECT 89.180 169.750 89.470 169.795 ;
        RECT 84.540 169.610 89.470 169.750 ;
        RECT 40.870 169.550 41.190 169.610 ;
        RECT 84.540 169.565 84.830 169.610 ;
        RECT 87.320 169.565 87.610 169.610 ;
        RECT 89.180 169.565 89.470 169.610 ;
        RECT 89.630 169.750 89.950 169.810 ;
        RECT 89.630 169.610 93.080 169.750 ;
        RECT 89.630 169.550 89.950 169.610 ;
        RECT 77.225 169.410 77.515 169.455 ;
        RECT 79.970 169.410 80.290 169.470 ;
        RECT 77.225 169.270 80.290 169.410 ;
        RECT 77.225 169.225 77.515 169.270 ;
        RECT 79.970 169.210 80.290 169.270 ;
        RECT 81.900 169.270 91.700 169.410 ;
        RECT 27.085 169.070 27.375 169.115 ;
        RECT 30.290 169.070 30.610 169.130 ;
        RECT 33.525 169.070 33.815 169.115 ;
        RECT 35.810 169.070 36.130 169.130 ;
        RECT 27.085 168.930 36.130 169.070 ;
        RECT 27.085 168.885 27.375 168.930 ;
        RECT 30.290 168.870 30.610 168.930 ;
        RECT 33.525 168.885 33.815 168.930 ;
        RECT 35.810 168.870 36.130 168.930 ;
        RECT 44.090 168.870 44.410 169.130 ;
        RECT 69.865 169.070 70.155 169.115 ;
        RECT 70.310 169.070 70.630 169.130 ;
        RECT 71.705 169.070 71.995 169.115 ;
        RECT 69.865 168.930 71.995 169.070 ;
        RECT 69.865 168.885 70.155 168.930 ;
        RECT 70.310 168.870 70.630 168.930 ;
        RECT 71.705 168.885 71.995 168.930 ;
        RECT 80.675 168.730 80.965 168.775 ;
        RECT 81.900 168.730 82.040 169.270 ;
        RECT 84.540 169.070 84.830 169.115 ;
        RECT 84.540 168.930 87.075 169.070 ;
        RECT 84.540 168.885 84.830 168.930 ;
        RECT 77.760 168.590 82.040 168.730 ;
        RECT 82.680 168.730 82.970 168.775 ;
        RECT 84.110 168.730 84.430 168.790 ;
        RECT 86.860 168.775 87.075 168.930 ;
        RECT 87.790 168.870 88.110 169.130 ;
        RECT 89.645 169.070 89.935 169.115 ;
        RECT 91.010 169.070 91.330 169.130 ;
        RECT 89.645 168.930 91.330 169.070 ;
        RECT 91.560 169.070 91.700 169.270 ;
        RECT 91.930 169.210 92.250 169.470 ;
        RECT 92.940 169.455 93.080 169.610 ;
        RECT 95.165 169.565 95.455 169.795 ;
        RECT 105.845 169.750 106.135 169.795 ;
        RECT 108.965 169.750 109.255 169.795 ;
        RECT 110.855 169.750 111.145 169.795 ;
        RECT 105.845 169.610 111.145 169.750 ;
        RECT 105.845 169.565 106.135 169.610 ;
        RECT 108.965 169.565 109.255 169.610 ;
        RECT 110.855 169.565 111.145 169.610 ;
        RECT 92.865 169.225 93.155 169.455 ;
        RECT 93.325 169.070 93.615 169.115 ;
        RECT 91.560 168.930 93.615 169.070 ;
        RECT 95.240 169.070 95.380 169.565 ;
        RECT 109.870 169.410 110.190 169.470 ;
        RECT 110.345 169.410 110.635 169.455 ;
        RECT 109.870 169.270 110.635 169.410 ;
        RECT 109.870 169.210 110.190 169.270 ;
        RECT 110.345 169.225 110.635 169.270 ;
        RECT 112.630 169.410 112.950 169.470 ;
        RECT 115.405 169.410 115.695 169.455 ;
        RECT 112.630 169.270 115.695 169.410 ;
        RECT 112.630 169.210 112.950 169.270 ;
        RECT 115.405 169.225 115.695 169.270 ;
        RECT 117.230 169.410 117.550 169.470 ;
        RECT 119.545 169.410 119.835 169.455 ;
        RECT 117.230 169.270 119.835 169.410 ;
        RECT 117.230 169.210 117.550 169.270 ;
        RECT 119.545 169.225 119.835 169.270 ;
        RECT 96.085 169.070 96.375 169.115 ;
        RECT 95.240 168.930 96.375 169.070 ;
        RECT 89.645 168.885 89.935 168.930 ;
        RECT 91.010 168.870 91.330 168.930 ;
        RECT 93.325 168.885 93.615 168.930 ;
        RECT 96.085 168.885 96.375 168.930 ;
        RECT 104.765 168.775 105.055 169.090 ;
        RECT 105.845 169.070 106.135 169.115 ;
        RECT 109.425 169.070 109.715 169.115 ;
        RECT 111.260 169.070 111.550 169.115 ;
        RECT 105.845 168.930 111.550 169.070 ;
        RECT 105.845 168.885 106.135 168.930 ;
        RECT 109.425 168.885 109.715 168.930 ;
        RECT 111.260 168.885 111.550 168.930 ;
        RECT 111.710 168.870 112.030 169.130 ;
        RECT 114.470 168.870 114.790 169.130 ;
        RECT 114.945 169.070 115.235 169.115 ;
        RECT 116.785 169.070 117.075 169.115 ;
        RECT 114.945 168.930 117.075 169.070 ;
        RECT 114.945 168.885 115.235 168.930 ;
        RECT 116.785 168.885 117.075 168.930 ;
        RECT 120.465 168.885 120.755 169.115 ;
        RECT 122.765 169.070 123.055 169.115 ;
        RECT 127.810 169.070 128.130 169.130 ;
        RECT 122.765 168.930 128.130 169.070 ;
        RECT 122.765 168.885 123.055 168.930 ;
        RECT 85.940 168.730 86.230 168.775 ;
        RECT 82.680 168.590 86.230 168.730 ;
        RECT 27.545 168.390 27.835 168.435 ;
        RECT 29.830 168.390 30.150 168.450 ;
        RECT 27.545 168.250 30.150 168.390 ;
        RECT 27.545 168.205 27.835 168.250 ;
        RECT 29.830 168.190 30.150 168.250 ;
        RECT 33.065 168.390 33.355 168.435 ;
        RECT 33.970 168.390 34.290 168.450 ;
        RECT 33.065 168.250 34.290 168.390 ;
        RECT 33.065 168.205 33.355 168.250 ;
        RECT 33.970 168.190 34.290 168.250 ;
        RECT 36.730 168.190 37.050 168.450 ;
        RECT 76.290 168.390 76.610 168.450 ;
        RECT 77.760 168.435 77.900 168.590 ;
        RECT 80.675 168.545 80.965 168.590 ;
        RECT 82.680 168.545 82.970 168.590 ;
        RECT 84.110 168.530 84.430 168.590 ;
        RECT 85.940 168.545 86.230 168.590 ;
        RECT 86.860 168.730 87.150 168.775 ;
        RECT 88.720 168.730 89.010 168.775 ;
        RECT 86.860 168.590 89.010 168.730 ;
        RECT 86.860 168.545 87.150 168.590 ;
        RECT 88.720 168.545 89.010 168.590 ;
        RECT 104.465 168.730 105.055 168.775 ;
        RECT 107.110 168.730 107.430 168.790 ;
        RECT 107.705 168.730 108.355 168.775 ;
        RECT 104.465 168.590 108.355 168.730 ;
        RECT 104.465 168.545 104.755 168.590 ;
        RECT 107.110 168.530 107.430 168.590 ;
        RECT 107.705 168.545 108.355 168.590 ;
        RECT 110.330 168.730 110.650 168.790 ;
        RECT 120.540 168.730 120.680 168.885 ;
        RECT 127.810 168.870 128.130 168.930 ;
        RECT 110.330 168.590 120.680 168.730 ;
        RECT 110.330 168.530 110.650 168.590 ;
        RECT 77.685 168.390 77.975 168.435 ;
        RECT 76.290 168.250 77.975 168.390 ;
        RECT 76.290 168.190 76.610 168.250 ;
        RECT 77.685 168.205 77.975 168.250 ;
        RECT 78.145 168.390 78.435 168.435 ;
        RECT 79.050 168.390 79.370 168.450 ;
        RECT 78.145 168.250 79.370 168.390 ;
        RECT 78.145 168.205 78.435 168.250 ;
        RECT 79.050 168.190 79.370 168.250 ;
        RECT 79.985 168.390 80.275 168.435 ;
        RECT 83.190 168.390 83.510 168.450 ;
        RECT 79.985 168.250 83.510 168.390 ;
        RECT 79.985 168.205 80.275 168.250 ;
        RECT 83.190 168.190 83.510 168.250 ;
        RECT 102.510 168.390 102.830 168.450 ;
        RECT 102.985 168.390 103.275 168.435 ;
        RECT 102.510 168.250 103.275 168.390 ;
        RECT 102.510 168.190 102.830 168.250 ;
        RECT 102.985 168.205 103.275 168.250 ;
        RECT 110.790 168.390 111.110 168.450 ;
        RECT 112.645 168.390 112.935 168.435 ;
        RECT 110.790 168.250 112.935 168.390 ;
        RECT 110.790 168.190 111.110 168.250 ;
        RECT 112.645 168.205 112.935 168.250 ;
        RECT 113.090 168.390 113.410 168.450 ;
        RECT 122.305 168.390 122.595 168.435 ;
        RECT 113.090 168.250 122.595 168.390 ;
        RECT 113.090 168.190 113.410 168.250 ;
        RECT 122.305 168.205 122.595 168.250 ;
        RECT 14.580 167.570 127.740 168.050 ;
        RECT 70.310 167.370 70.630 167.430 ;
        RECT 48.320 167.230 53.060 167.370 ;
        RECT 24.770 166.830 25.090 167.090 ;
        RECT 27.065 167.030 27.715 167.075 ;
        RECT 29.830 167.030 30.150 167.090 ;
        RECT 30.665 167.030 30.955 167.075 ;
        RECT 27.065 166.890 30.955 167.030 ;
        RECT 27.065 166.845 27.715 166.890 ;
        RECT 29.830 166.830 30.150 166.890 ;
        RECT 30.365 166.845 30.955 166.890 ;
        RECT 35.810 167.030 36.130 167.090 ;
        RECT 48.320 167.030 48.460 167.230 ;
        RECT 35.810 166.890 48.460 167.030 ;
        RECT 48.805 167.030 49.095 167.075 ;
        RECT 50.990 167.030 51.310 167.090 ;
        RECT 52.045 167.030 52.695 167.075 ;
        RECT 48.805 166.890 52.695 167.030 ;
        RECT 52.920 167.030 53.060 167.230 ;
        RECT 70.310 167.230 73.760 167.370 ;
        RECT 70.310 167.170 70.630 167.230 ;
        RECT 53.290 167.030 53.610 167.090 ;
        RECT 73.085 167.030 73.375 167.075 ;
        RECT 52.920 166.890 59.500 167.030 ;
        RECT 23.870 166.690 24.160 166.735 ;
        RECT 25.705 166.690 25.995 166.735 ;
        RECT 29.285 166.690 29.575 166.735 ;
        RECT 23.870 166.550 29.575 166.690 ;
        RECT 23.870 166.505 24.160 166.550 ;
        RECT 25.705 166.505 25.995 166.550 ;
        RECT 29.285 166.505 29.575 166.550 ;
        RECT 30.365 166.530 30.655 166.845 ;
        RECT 35.810 166.830 36.130 166.890 ;
        RECT 33.525 166.690 33.815 166.735 ;
        RECT 34.430 166.690 34.750 166.750 ;
        RECT 33.525 166.550 34.750 166.690 ;
        RECT 33.525 166.505 33.815 166.550 ;
        RECT 34.430 166.490 34.750 166.550 ;
        RECT 36.285 166.690 36.575 166.735 ;
        RECT 36.730 166.690 37.050 166.750 ;
        RECT 37.740 166.735 37.880 166.890 ;
        RECT 48.805 166.845 49.395 166.890 ;
        RECT 36.285 166.550 37.050 166.690 ;
        RECT 36.285 166.505 36.575 166.550 ;
        RECT 36.730 166.490 37.050 166.550 ;
        RECT 37.665 166.505 37.955 166.735 ;
        RECT 45.560 166.550 48.920 166.690 ;
        RECT 23.405 166.350 23.695 166.395 ;
        RECT 27.070 166.350 27.390 166.410 ;
        RECT 23.405 166.210 27.390 166.350 ;
        RECT 23.405 166.165 23.695 166.210 ;
        RECT 27.070 166.150 27.390 166.210 ;
        RECT 32.145 166.350 32.435 166.395 ;
        RECT 39.505 166.350 39.795 166.395 ;
        RECT 43.170 166.350 43.490 166.410 ;
        RECT 32.145 166.210 43.490 166.350 ;
        RECT 32.145 166.165 32.435 166.210 ;
        RECT 39.505 166.165 39.795 166.210 ;
        RECT 43.170 166.150 43.490 166.210 ;
        RECT 24.275 166.010 24.565 166.055 ;
        RECT 26.165 166.010 26.455 166.055 ;
        RECT 29.285 166.010 29.575 166.055 ;
        RECT 24.275 165.870 29.575 166.010 ;
        RECT 24.275 165.825 24.565 165.870 ;
        RECT 26.165 165.825 26.455 165.870 ;
        RECT 29.285 165.825 29.575 165.870 ;
        RECT 29.830 166.010 30.150 166.070 ;
        RECT 42.265 166.010 42.555 166.055 ;
        RECT 45.560 166.010 45.700 166.550 ;
        RECT 45.945 166.350 46.235 166.395 ;
        RECT 48.780 166.350 48.920 166.550 ;
        RECT 49.105 166.530 49.395 166.845 ;
        RECT 50.990 166.830 51.310 166.890 ;
        RECT 52.045 166.845 52.695 166.890 ;
        RECT 53.290 166.830 53.610 166.890 ;
        RECT 59.360 166.735 59.500 166.890 ;
        RECT 68.560 166.890 73.375 167.030 ;
        RECT 68.560 166.750 68.700 166.890 ;
        RECT 73.085 166.845 73.375 166.890 ;
        RECT 50.185 166.690 50.475 166.735 ;
        RECT 53.765 166.690 54.055 166.735 ;
        RECT 55.600 166.690 55.890 166.735 ;
        RECT 50.185 166.550 55.890 166.690 ;
        RECT 50.185 166.505 50.475 166.550 ;
        RECT 53.765 166.505 54.055 166.550 ;
        RECT 55.600 166.505 55.890 166.550 ;
        RECT 59.285 166.690 59.575 166.735 ;
        RECT 61.125 166.690 61.415 166.735 ;
        RECT 59.285 166.550 61.415 166.690 ;
        RECT 59.285 166.505 59.575 166.550 ;
        RECT 61.125 166.505 61.415 166.550 ;
        RECT 61.570 166.690 61.890 166.750 ;
        RECT 62.505 166.690 62.795 166.735 ;
        RECT 67.105 166.690 67.395 166.735 ;
        RECT 61.570 166.550 67.395 166.690 ;
        RECT 61.570 166.490 61.890 166.550 ;
        RECT 62.505 166.505 62.795 166.550 ;
        RECT 67.105 166.505 67.395 166.550 ;
        RECT 68.470 166.490 68.790 166.750 ;
        RECT 70.770 166.490 71.090 166.750 ;
        RECT 72.625 166.690 72.915 166.735 ;
        RECT 73.620 166.690 73.760 167.230 ;
        RECT 110.330 167.170 110.650 167.430 ;
        RECT 77.620 167.030 77.910 167.075 ;
        RECT 80.880 167.030 81.170 167.075 ;
        RECT 77.620 166.890 81.170 167.030 ;
        RECT 77.620 166.845 77.910 166.890 ;
        RECT 72.625 166.550 73.760 166.690 ;
        RECT 72.625 166.505 72.915 166.550 ;
        RECT 54.210 166.350 54.530 166.410 ;
        RECT 45.945 166.210 47.540 166.350 ;
        RECT 48.780 166.210 54.530 166.350 ;
        RECT 45.945 166.165 46.235 166.210 ;
        RECT 29.830 165.870 45.700 166.010 ;
        RECT 29.830 165.810 30.150 165.870 ;
        RECT 42.265 165.825 42.555 165.870 ;
        RECT 28.450 165.670 28.770 165.730 ;
        RECT 32.605 165.670 32.895 165.715 ;
        RECT 28.450 165.530 32.895 165.670 ;
        RECT 28.450 165.470 28.770 165.530 ;
        RECT 32.605 165.485 32.895 165.530 ;
        RECT 38.110 165.470 38.430 165.730 ;
        RECT 42.710 165.470 43.030 165.730 ;
        RECT 47.400 165.715 47.540 166.210 ;
        RECT 54.210 166.150 54.530 166.210 ;
        RECT 54.670 166.150 54.990 166.410 ;
        RECT 56.065 166.350 56.355 166.395 ;
        RECT 57.430 166.350 57.750 166.410 ;
        RECT 63.870 166.350 64.190 166.410 ;
        RECT 56.065 166.210 64.190 166.350 ;
        RECT 56.065 166.165 56.355 166.210 ;
        RECT 57.430 166.150 57.750 166.210 ;
        RECT 63.870 166.150 64.190 166.210 ;
        RECT 66.630 166.350 66.950 166.410 ;
        RECT 71.245 166.350 71.535 166.395 ;
        RECT 66.630 166.210 71.535 166.350 ;
        RECT 66.630 166.150 66.950 166.210 ;
        RECT 71.245 166.165 71.535 166.210 ;
        RECT 72.165 166.350 72.455 166.395 ;
        RECT 73.990 166.350 74.310 166.410 ;
        RECT 74.910 166.350 75.230 166.410 ;
        RECT 72.165 166.210 75.230 166.350 ;
        RECT 79.140 166.350 79.280 166.890 ;
        RECT 80.880 166.845 81.170 166.890 ;
        RECT 81.800 167.030 82.090 167.075 ;
        RECT 83.660 167.030 83.950 167.075 ;
        RECT 81.800 166.890 83.950 167.030 ;
        RECT 81.800 166.845 82.090 166.890 ;
        RECT 83.660 166.845 83.950 166.890 ;
        RECT 84.110 167.030 84.430 167.090 ;
        RECT 86.885 167.030 87.175 167.075 ;
        RECT 84.110 166.890 87.175 167.030 ;
        RECT 79.480 166.690 79.770 166.735 ;
        RECT 81.800 166.690 82.015 166.845 ;
        RECT 84.110 166.830 84.430 166.890 ;
        RECT 86.885 166.845 87.175 166.890 ;
        RECT 99.700 167.030 99.990 167.075 ;
        RECT 100.210 167.030 100.530 167.090 ;
        RECT 102.960 167.030 103.250 167.075 ;
        RECT 99.700 166.890 103.250 167.030 ;
        RECT 99.700 166.845 99.990 166.890 ;
        RECT 100.210 166.830 100.530 166.890 ;
        RECT 102.960 166.845 103.250 166.890 ;
        RECT 103.880 167.030 104.170 167.075 ;
        RECT 105.740 167.030 106.030 167.075 ;
        RECT 103.880 166.890 106.030 167.030 ;
        RECT 103.880 166.845 104.170 166.890 ;
        RECT 105.740 166.845 106.030 166.890 ;
        RECT 117.345 167.030 117.635 167.075 ;
        RECT 119.530 167.030 119.850 167.090 ;
        RECT 120.585 167.030 121.235 167.075 ;
        RECT 117.345 166.890 121.235 167.030 ;
        RECT 117.345 166.845 117.935 166.890 ;
        RECT 85.505 166.690 85.795 166.735 ;
        RECT 79.480 166.550 82.015 166.690 ;
        RECT 82.360 166.550 85.795 166.690 ;
        RECT 79.480 166.505 79.770 166.550 ;
        RECT 82.360 166.350 82.500 166.550 ;
        RECT 85.505 166.505 85.795 166.550 ;
        RECT 85.965 166.690 86.255 166.735 ;
        RECT 87.345 166.690 87.635 166.735 ;
        RECT 88.710 166.690 89.030 166.750 ;
        RECT 85.965 166.550 89.030 166.690 ;
        RECT 85.965 166.505 86.255 166.550 ;
        RECT 87.345 166.505 87.635 166.550 ;
        RECT 88.710 166.490 89.030 166.550 ;
        RECT 95.165 166.505 95.455 166.735 ;
        RECT 101.560 166.690 101.850 166.735 ;
        RECT 103.880 166.690 104.095 166.845 ;
        RECT 101.560 166.550 104.095 166.690 ;
        RECT 107.585 166.690 107.875 166.735 ;
        RECT 110.790 166.690 111.110 166.750 ;
        RECT 107.585 166.550 111.110 166.690 ;
        RECT 101.560 166.505 101.850 166.550 ;
        RECT 107.585 166.505 107.875 166.550 ;
        RECT 79.140 166.210 82.500 166.350 ;
        RECT 72.165 166.165 72.455 166.210 ;
        RECT 73.990 166.150 74.310 166.210 ;
        RECT 74.910 166.150 75.230 166.210 ;
        RECT 82.730 166.150 83.050 166.410 ;
        RECT 84.585 166.350 84.875 166.395 ;
        RECT 91.010 166.350 91.330 166.410 ;
        RECT 84.585 166.210 91.330 166.350 ;
        RECT 84.585 166.165 84.875 166.210 ;
        RECT 91.010 166.150 91.330 166.210 ;
        RECT 91.930 166.350 92.250 166.410 ;
        RECT 93.770 166.350 94.090 166.410 ;
        RECT 91.930 166.210 94.090 166.350 ;
        RECT 91.930 166.150 92.250 166.210 ;
        RECT 93.770 166.150 94.090 166.210 ;
        RECT 94.690 166.150 95.010 166.410 ;
        RECT 95.240 166.350 95.380 166.505 ;
        RECT 110.790 166.490 111.110 166.550 ;
        RECT 111.265 166.690 111.555 166.735 ;
        RECT 112.170 166.690 112.490 166.750 ;
        RECT 111.265 166.550 112.490 166.690 ;
        RECT 111.265 166.505 111.555 166.550 ;
        RECT 112.170 166.490 112.490 166.550 ;
        RECT 117.645 166.530 117.935 166.845 ;
        RECT 119.530 166.830 119.850 166.890 ;
        RECT 120.585 166.845 121.235 166.890 ;
        RECT 118.725 166.690 119.015 166.735 ;
        RECT 122.305 166.690 122.595 166.735 ;
        RECT 124.140 166.690 124.430 166.735 ;
        RECT 118.725 166.550 124.430 166.690 ;
        RECT 118.725 166.505 119.015 166.550 ;
        RECT 122.305 166.505 122.595 166.550 ;
        RECT 124.140 166.505 124.430 166.550 ;
        RECT 124.590 166.490 124.910 166.750 ;
        RECT 97.695 166.350 97.985 166.395 ;
        RECT 98.370 166.350 98.690 166.410 ;
        RECT 95.240 166.210 98.690 166.350 ;
        RECT 97.695 166.165 97.985 166.210 ;
        RECT 98.370 166.150 98.690 166.210 ;
        RECT 104.810 166.150 105.130 166.410 ;
        RECT 105.730 166.350 106.050 166.410 ;
        RECT 106.665 166.350 106.955 166.395 ;
        RECT 111.710 166.350 112.030 166.410 ;
        RECT 124.680 166.350 124.820 166.490 ;
        RECT 105.730 166.210 124.820 166.350 ;
        RECT 105.730 166.150 106.050 166.210 ;
        RECT 106.665 166.165 106.955 166.210 ;
        RECT 111.710 166.150 112.030 166.210 ;
        RECT 50.185 166.010 50.475 166.055 ;
        RECT 53.305 166.010 53.595 166.055 ;
        RECT 55.195 166.010 55.485 166.055 ;
        RECT 50.185 165.870 55.485 166.010 ;
        RECT 50.185 165.825 50.475 165.870 ;
        RECT 53.305 165.825 53.595 165.870 ;
        RECT 55.195 165.825 55.485 165.870 ;
        RECT 69.865 166.010 70.155 166.055 ;
        RECT 78.590 166.010 78.910 166.070 ;
        RECT 69.865 165.870 78.910 166.010 ;
        RECT 69.865 165.825 70.155 165.870 ;
        RECT 78.590 165.810 78.910 165.870 ;
        RECT 79.480 166.010 79.770 166.055 ;
        RECT 82.260 166.010 82.550 166.055 ;
        RECT 84.120 166.010 84.410 166.055 ;
        RECT 79.480 165.870 84.410 166.010 ;
        RECT 79.480 165.825 79.770 165.870 ;
        RECT 82.260 165.825 82.550 165.870 ;
        RECT 84.120 165.825 84.410 165.870 ;
        RECT 101.560 166.010 101.850 166.055 ;
        RECT 104.340 166.010 104.630 166.055 ;
        RECT 106.200 166.010 106.490 166.055 ;
        RECT 101.560 165.870 106.490 166.010 ;
        RECT 101.560 165.825 101.850 165.870 ;
        RECT 104.340 165.825 104.630 165.870 ;
        RECT 106.200 165.825 106.490 165.870 ;
        RECT 108.950 166.010 109.270 166.070 ;
        RECT 110.790 166.010 111.110 166.070 ;
        RECT 108.950 165.870 111.110 166.010 ;
        RECT 108.950 165.810 109.270 165.870 ;
        RECT 110.790 165.810 111.110 165.870 ;
        RECT 112.170 166.010 112.490 166.070 ;
        RECT 115.865 166.010 116.155 166.055 ;
        RECT 112.170 165.870 116.155 166.010 ;
        RECT 112.170 165.810 112.490 165.870 ;
        RECT 115.865 165.825 116.155 165.870 ;
        RECT 118.725 166.010 119.015 166.055 ;
        RECT 121.845 166.010 122.135 166.055 ;
        RECT 123.735 166.010 124.025 166.055 ;
        RECT 118.725 165.870 124.025 166.010 ;
        RECT 118.725 165.825 119.015 165.870 ;
        RECT 121.845 165.825 122.135 165.870 ;
        RECT 123.735 165.825 124.025 165.870 ;
        RECT 47.325 165.670 47.615 165.715 ;
        RECT 49.610 165.670 49.930 165.730 ;
        RECT 47.325 165.530 49.930 165.670 ;
        RECT 47.325 165.485 47.615 165.530 ;
        RECT 49.610 165.470 49.930 165.530 ;
        RECT 58.810 165.470 59.130 165.730 ;
        RECT 66.645 165.670 66.935 165.715 ;
        RECT 68.930 165.670 69.250 165.730 ;
        RECT 66.645 165.530 69.250 165.670 ;
        RECT 66.645 165.485 66.935 165.530 ;
        RECT 68.930 165.470 69.250 165.530 ;
        RECT 73.070 165.670 73.390 165.730 ;
        RECT 75.615 165.670 75.905 165.715 ;
        RECT 73.070 165.530 75.905 165.670 ;
        RECT 78.680 165.670 78.820 165.810 ;
        RECT 79.970 165.670 80.290 165.730 ;
        RECT 91.930 165.670 92.250 165.730 ;
        RECT 78.680 165.530 92.250 165.670 ;
        RECT 73.070 165.470 73.390 165.530 ;
        RECT 75.615 165.485 75.905 165.530 ;
        RECT 79.970 165.470 80.290 165.530 ;
        RECT 91.930 165.470 92.250 165.530 ;
        RECT 96.530 165.670 96.850 165.730 ;
        RECT 97.005 165.670 97.295 165.715 ;
        RECT 96.530 165.530 97.295 165.670 ;
        RECT 96.530 165.470 96.850 165.530 ;
        RECT 97.005 165.485 97.295 165.530 ;
        RECT 114.010 165.470 114.330 165.730 ;
        RECT 121.370 165.670 121.690 165.730 ;
        RECT 123.290 165.670 123.580 165.715 ;
        RECT 121.370 165.530 123.580 165.670 ;
        RECT 121.370 165.470 121.690 165.530 ;
        RECT 123.290 165.485 123.580 165.530 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 14.580 164.850 127.740 165.330 ;
        RECT 24.770 164.650 25.090 164.710 ;
        RECT 25.705 164.650 25.995 164.695 ;
        RECT 24.770 164.510 25.995 164.650 ;
        RECT 24.770 164.450 25.090 164.510 ;
        RECT 25.705 164.465 25.995 164.510 ;
        RECT 50.990 164.450 51.310 164.710 ;
        RECT 54.670 164.450 54.990 164.710 ;
        RECT 61.570 164.650 61.890 164.710 ;
        RECT 82.730 164.650 83.050 164.710 ;
        RECT 83.205 164.650 83.495 164.695 ;
        RECT 61.570 164.510 71.230 164.650 ;
        RECT 61.570 164.450 61.890 164.510 ;
        RECT 27.955 164.310 28.245 164.355 ;
        RECT 29.845 164.310 30.135 164.355 ;
        RECT 32.965 164.310 33.255 164.355 ;
        RECT 27.955 164.170 33.255 164.310 ;
        RECT 27.955 164.125 28.245 164.170 ;
        RECT 29.845 164.125 30.135 164.170 ;
        RECT 32.965 164.125 33.255 164.170 ;
        RECT 39.145 164.310 39.435 164.355 ;
        RECT 42.265 164.310 42.555 164.355 ;
        RECT 44.155 164.310 44.445 164.355 ;
        RECT 57.430 164.310 57.750 164.370 ;
        RECT 39.145 164.170 44.445 164.310 ;
        RECT 39.145 164.125 39.435 164.170 ;
        RECT 42.265 164.125 42.555 164.170 ;
        RECT 44.155 164.125 44.445 164.170 ;
        RECT 45.100 164.170 57.750 164.310 ;
        RECT 28.450 163.770 28.770 164.030 ;
        RECT 28.910 163.970 29.230 164.030 ;
        RECT 36.730 163.970 37.050 164.030 ;
        RECT 45.100 164.015 45.240 164.170 ;
        RECT 57.430 164.110 57.750 164.170 ;
        RECT 58.005 164.310 58.295 164.355 ;
        RECT 61.125 164.310 61.415 164.355 ;
        RECT 63.015 164.310 63.305 164.355 ;
        RECT 58.005 164.170 63.305 164.310 ;
        RECT 58.005 164.125 58.295 164.170 ;
        RECT 61.125 164.125 61.415 164.170 ;
        RECT 63.015 164.125 63.305 164.170 ;
        RECT 45.025 163.970 45.315 164.015 ;
        RECT 28.910 163.830 45.315 163.970 ;
        RECT 28.910 163.770 29.230 163.830 ;
        RECT 36.730 163.770 37.050 163.830 ;
        RECT 45.025 163.785 45.315 163.830 ;
        RECT 49.625 163.970 49.915 164.015 ;
        RECT 60.650 163.970 60.970 164.030 ;
        RECT 49.625 163.830 53.980 163.970 ;
        RECT 49.625 163.785 49.915 163.830 ;
        RECT 26.610 163.430 26.930 163.690 ;
        RECT 27.070 163.430 27.390 163.690 ;
        RECT 27.550 163.630 27.840 163.675 ;
        RECT 29.385 163.630 29.675 163.675 ;
        RECT 32.965 163.630 33.255 163.675 ;
        RECT 27.550 163.490 33.255 163.630 ;
        RECT 27.550 163.445 27.840 163.490 ;
        RECT 29.385 163.445 29.675 163.490 ;
        RECT 32.965 163.445 33.255 163.490 ;
        RECT 33.970 163.650 34.290 163.690 ;
        RECT 38.110 163.650 38.430 163.690 ;
        RECT 33.970 163.430 34.335 163.650 ;
        RECT 27.160 163.290 27.300 163.430 ;
        RECT 28.910 163.290 29.230 163.350 ;
        RECT 34.045 163.335 34.335 163.430 ;
        RECT 38.065 163.430 38.430 163.650 ;
        RECT 39.145 163.630 39.435 163.675 ;
        RECT 42.725 163.630 43.015 163.675 ;
        RECT 44.560 163.630 44.850 163.675 ;
        RECT 39.145 163.490 44.850 163.630 ;
        RECT 39.145 163.445 39.435 163.490 ;
        RECT 42.725 163.445 43.015 163.490 ;
        RECT 44.560 163.445 44.850 163.490 ;
        RECT 46.865 163.630 47.155 163.675 ;
        RECT 49.150 163.630 49.470 163.690 ;
        RECT 46.865 163.490 49.470 163.630 ;
        RECT 46.865 163.445 47.155 163.490 ;
        RECT 49.150 163.430 49.470 163.490 ;
        RECT 51.465 163.630 51.755 163.675 ;
        RECT 53.290 163.630 53.610 163.690 ;
        RECT 53.840 163.675 53.980 163.830 ;
        RECT 60.650 163.830 65.480 163.970 ;
        RECT 60.650 163.770 60.970 163.830 ;
        RECT 51.465 163.490 53.610 163.630 ;
        RECT 51.465 163.445 51.755 163.490 ;
        RECT 53.290 163.430 53.610 163.490 ;
        RECT 53.765 163.445 54.055 163.675 ;
        RECT 38.065 163.335 38.355 163.430 ;
        RECT 27.160 163.150 29.230 163.290 ;
        RECT 28.910 163.090 29.230 163.150 ;
        RECT 30.745 163.290 31.395 163.335 ;
        RECT 34.045 163.290 34.635 163.335 ;
        RECT 30.745 163.150 34.635 163.290 ;
        RECT 30.745 163.105 31.395 163.150 ;
        RECT 34.345 163.105 34.635 163.150 ;
        RECT 37.765 163.290 38.355 163.335 ;
        RECT 41.005 163.290 41.655 163.335 ;
        RECT 37.765 163.150 41.655 163.290 ;
        RECT 37.765 163.105 38.055 163.150 ;
        RECT 41.005 163.105 41.655 163.150 ;
        RECT 43.645 163.290 43.935 163.335 ;
        RECT 46.390 163.290 46.710 163.350 ;
        RECT 56.925 163.335 57.215 163.650 ;
        RECT 58.005 163.630 58.295 163.675 ;
        RECT 61.585 163.630 61.875 163.675 ;
        RECT 63.420 163.630 63.710 163.675 ;
        RECT 58.005 163.490 63.710 163.630 ;
        RECT 58.005 163.445 58.295 163.490 ;
        RECT 61.585 163.445 61.875 163.490 ;
        RECT 63.420 163.445 63.710 163.490 ;
        RECT 63.870 163.430 64.190 163.690 ;
        RECT 43.645 163.150 46.710 163.290 ;
        RECT 43.645 163.105 43.935 163.150 ;
        RECT 46.390 163.090 46.710 163.150 ;
        RECT 56.625 163.290 57.215 163.335 ;
        RECT 58.810 163.290 59.130 163.350 ;
        RECT 59.865 163.290 60.515 163.335 ;
        RECT 56.625 163.150 60.515 163.290 ;
        RECT 56.625 163.105 56.915 163.150 ;
        RECT 58.810 163.090 59.130 163.150 ;
        RECT 59.865 163.105 60.515 163.150 ;
        RECT 62.490 163.090 62.810 163.350 ;
        RECT 65.340 163.335 65.480 163.830 ;
        RECT 65.800 163.630 65.940 164.510 ;
        RECT 71.090 164.310 71.230 164.510 ;
        RECT 82.730 164.510 83.495 164.650 ;
        RECT 82.730 164.450 83.050 164.510 ;
        RECT 83.205 164.465 83.495 164.510 ;
        RECT 86.425 164.650 86.715 164.695 ;
        RECT 87.790 164.650 88.110 164.710 ;
        RECT 113.090 164.650 113.410 164.710 ;
        RECT 86.425 164.510 88.110 164.650 ;
        RECT 86.425 164.465 86.715 164.510 ;
        RECT 87.790 164.450 88.110 164.510 ;
        RECT 105.820 164.510 113.410 164.650 ;
        RECT 105.820 164.310 105.960 164.510 ;
        RECT 113.090 164.450 113.410 164.510 ;
        RECT 71.090 164.170 105.960 164.310 ;
        RECT 106.665 164.310 106.955 164.355 ;
        RECT 108.950 164.310 109.270 164.370 ;
        RECT 106.665 164.170 109.270 164.310 ;
        RECT 106.665 164.125 106.955 164.170 ;
        RECT 108.950 164.110 109.270 164.170 ;
        RECT 116.425 164.310 116.715 164.355 ;
        RECT 119.545 164.310 119.835 164.355 ;
        RECT 121.435 164.310 121.725 164.355 ;
        RECT 116.425 164.170 121.725 164.310 ;
        RECT 116.425 164.125 116.715 164.170 ;
        RECT 119.545 164.125 119.835 164.170 ;
        RECT 121.435 164.125 121.725 164.170 ;
        RECT 78.590 163.770 78.910 164.030 ;
        RECT 93.770 163.970 94.090 164.030 ;
        RECT 102.525 163.970 102.815 164.015 ;
        RECT 109.425 163.970 109.715 164.015 ;
        RECT 93.770 163.830 109.715 163.970 ;
        RECT 93.770 163.770 94.090 163.830 ;
        RECT 102.525 163.785 102.815 163.830 ;
        RECT 109.425 163.785 109.715 163.830 ;
        RECT 110.330 163.970 110.650 164.030 ;
        RECT 113.565 163.970 113.855 164.015 ;
        RECT 110.330 163.830 113.855 163.970 ;
        RECT 66.645 163.630 66.935 163.675 ;
        RECT 65.800 163.490 66.935 163.630 ;
        RECT 66.645 163.445 66.935 163.490 ;
        RECT 68.470 163.630 68.790 163.690 ;
        RECT 68.945 163.630 69.235 163.675 ;
        RECT 68.470 163.490 69.235 163.630 ;
        RECT 68.470 163.430 68.790 163.490 ;
        RECT 68.945 163.445 69.235 163.490 ;
        RECT 73.070 163.630 73.390 163.690 ;
        RECT 79.525 163.630 79.815 163.675 ;
        RECT 82.285 163.630 82.575 163.675 ;
        RECT 73.070 163.490 79.815 163.630 ;
        RECT 73.070 163.430 73.390 163.490 ;
        RECT 79.140 163.350 79.280 163.490 ;
        RECT 79.525 163.445 79.815 163.490 ;
        RECT 81.900 163.490 82.575 163.630 ;
        RECT 65.265 163.290 65.555 163.335 ;
        RECT 75.370 163.290 75.690 163.350 ;
        RECT 65.265 163.150 75.690 163.290 ;
        RECT 65.265 163.105 65.555 163.150 ;
        RECT 75.370 163.090 75.690 163.150 ;
        RECT 79.050 163.090 79.370 163.350 ;
        RECT 35.810 162.750 36.130 163.010 ;
        RECT 36.270 162.750 36.590 163.010 ;
        RECT 52.830 162.950 53.150 163.010 ;
        RECT 55.145 162.950 55.435 162.995 ;
        RECT 52.830 162.810 55.435 162.950 ;
        RECT 52.830 162.750 53.150 162.810 ;
        RECT 55.145 162.765 55.435 162.810 ;
        RECT 67.090 162.950 67.410 163.010 ;
        RECT 67.565 162.950 67.855 162.995 ;
        RECT 67.090 162.810 67.855 162.950 ;
        RECT 67.090 162.750 67.410 162.810 ;
        RECT 67.565 162.765 67.855 162.810 ;
        RECT 79.985 162.950 80.275 162.995 ;
        RECT 80.890 162.950 81.210 163.010 ;
        RECT 81.900 162.995 82.040 163.490 ;
        RECT 82.285 163.445 82.575 163.490 ;
        RECT 83.190 163.630 83.510 163.690 ;
        RECT 85.505 163.630 85.795 163.675 ;
        RECT 83.190 163.490 85.795 163.630 ;
        RECT 83.190 163.430 83.510 163.490 ;
        RECT 85.505 163.445 85.795 163.490 ;
        RECT 101.130 163.430 101.450 163.690 ;
        RECT 109.500 163.630 109.640 163.785 ;
        RECT 110.330 163.770 110.650 163.830 ;
        RECT 113.565 163.785 113.855 163.830 ;
        RECT 122.305 163.970 122.595 164.015 ;
        RECT 124.590 163.970 124.910 164.030 ;
        RECT 122.305 163.830 124.910 163.970 ;
        RECT 122.305 163.785 122.595 163.830 ;
        RECT 124.590 163.770 124.910 163.830 ;
        RECT 112.630 163.630 112.950 163.690 ;
        RECT 109.500 163.490 112.950 163.630 ;
        RECT 112.630 163.430 112.950 163.490 ;
        RECT 113.090 163.430 113.410 163.690 ;
        RECT 98.370 163.290 98.690 163.350 ;
        RECT 103.445 163.290 103.735 163.335 ;
        RECT 98.370 163.150 103.735 163.290 ;
        RECT 98.370 163.090 98.690 163.150 ;
        RECT 103.445 163.105 103.735 163.150 ;
        RECT 103.905 163.290 104.195 163.335 ;
        RECT 106.190 163.290 106.510 163.350 ;
        RECT 108.965 163.290 109.255 163.335 ;
        RECT 103.905 163.150 109.255 163.290 ;
        RECT 103.905 163.105 104.195 163.150 ;
        RECT 106.190 163.090 106.510 163.150 ;
        RECT 108.965 163.105 109.255 163.150 ;
        RECT 111.710 163.090 112.030 163.350 ;
        RECT 113.550 163.290 113.870 163.350 ;
        RECT 115.345 163.335 115.635 163.650 ;
        RECT 116.425 163.630 116.715 163.675 ;
        RECT 120.005 163.630 120.295 163.675 ;
        RECT 121.840 163.630 122.130 163.675 ;
        RECT 116.425 163.490 122.130 163.630 ;
        RECT 116.425 163.445 116.715 163.490 ;
        RECT 120.005 163.445 120.295 163.490 ;
        RECT 121.840 163.445 122.130 163.490 ;
        RECT 123.670 163.430 123.990 163.690 ;
        RECT 115.045 163.290 115.635 163.335 ;
        RECT 118.285 163.290 118.935 163.335 ;
        RECT 113.550 163.150 118.935 163.290 ;
        RECT 113.550 163.090 113.870 163.150 ;
        RECT 115.045 163.105 115.335 163.150 ;
        RECT 118.285 163.105 118.935 163.150 ;
        RECT 120.925 163.105 121.215 163.335 ;
        RECT 79.985 162.810 81.210 162.950 ;
        RECT 79.985 162.765 80.275 162.810 ;
        RECT 80.890 162.750 81.210 162.810 ;
        RECT 81.825 162.765 82.115 162.995 ;
        RECT 91.010 162.950 91.330 163.010 ;
        RECT 94.705 162.950 94.995 162.995 ;
        RECT 97.450 162.950 97.770 163.010 ;
        RECT 91.010 162.810 97.770 162.950 ;
        RECT 91.010 162.750 91.330 162.810 ;
        RECT 94.705 162.765 94.995 162.810 ;
        RECT 97.450 162.750 97.770 162.810 ;
        RECT 105.270 162.950 105.590 163.010 ;
        RECT 105.745 162.950 106.035 162.995 ;
        RECT 105.270 162.810 106.035 162.950 ;
        RECT 105.270 162.750 105.590 162.810 ;
        RECT 105.745 162.765 106.035 162.810 ;
        RECT 108.505 162.950 108.795 162.995 ;
        RECT 109.870 162.950 110.190 163.010 ;
        RECT 108.505 162.810 110.190 162.950 ;
        RECT 121.000 162.950 121.140 163.105 ;
        RECT 122.765 162.950 123.055 162.995 ;
        RECT 121.000 162.810 123.055 162.950 ;
        RECT 108.505 162.765 108.795 162.810 ;
        RECT 109.870 162.750 110.190 162.810 ;
        RECT 122.765 162.765 123.055 162.810 ;
        RECT 14.580 162.130 127.740 162.610 ;
        RECT 26.610 161.930 26.930 161.990 ;
        RECT 27.545 161.930 27.835 161.975 ;
        RECT 26.610 161.790 27.835 161.930 ;
        RECT 26.610 161.730 26.930 161.790 ;
        RECT 27.545 161.745 27.835 161.790 ;
        RECT 29.830 161.730 30.150 161.990 ;
        RECT 33.065 161.930 33.355 161.975 ;
        RECT 34.430 161.930 34.750 161.990 ;
        RECT 33.065 161.790 34.750 161.930 ;
        RECT 33.065 161.745 33.355 161.790 ;
        RECT 34.430 161.730 34.750 161.790 ;
        RECT 42.710 161.930 43.030 161.990 ;
        RECT 45.485 161.930 45.775 161.975 ;
        RECT 42.710 161.790 45.775 161.930 ;
        RECT 42.710 161.730 43.030 161.790 ;
        RECT 45.485 161.745 45.775 161.790 ;
        RECT 46.390 161.930 46.710 161.990 ;
        RECT 47.785 161.930 48.075 161.975 ;
        RECT 46.390 161.790 48.075 161.930 ;
        RECT 46.390 161.730 46.710 161.790 ;
        RECT 47.785 161.745 48.075 161.790 ;
        RECT 49.150 161.730 49.470 161.990 ;
        RECT 49.610 161.730 49.930 161.990 ;
        RECT 54.210 161.930 54.530 161.990 ;
        RECT 55.145 161.930 55.435 161.975 ;
        RECT 54.210 161.790 55.435 161.930 ;
        RECT 54.210 161.730 54.530 161.790 ;
        RECT 55.145 161.745 55.435 161.790 ;
        RECT 56.985 161.745 57.275 161.975 ;
        RECT 60.665 161.930 60.955 161.975 ;
        RECT 62.490 161.930 62.810 161.990 ;
        RECT 60.665 161.790 62.810 161.930 ;
        RECT 60.665 161.745 60.955 161.790 ;
        RECT 18.790 161.590 19.110 161.650 ;
        RECT 20.120 161.590 20.410 161.635 ;
        RECT 23.380 161.590 23.670 161.635 ;
        RECT 18.790 161.450 23.670 161.590 ;
        RECT 18.790 161.390 19.110 161.450 ;
        RECT 20.120 161.405 20.410 161.450 ;
        RECT 23.380 161.405 23.670 161.450 ;
        RECT 24.300 161.590 24.590 161.635 ;
        RECT 26.160 161.590 26.450 161.635 ;
        RECT 24.300 161.450 26.450 161.590 ;
        RECT 24.300 161.405 24.590 161.450 ;
        RECT 26.160 161.405 26.450 161.450 ;
        RECT 29.385 161.405 29.675 161.635 ;
        RECT 31.210 161.590 31.530 161.650 ;
        RECT 34.905 161.590 35.195 161.635 ;
        RECT 31.210 161.450 35.195 161.590 ;
        RECT 21.980 161.250 22.270 161.295 ;
        RECT 24.300 161.250 24.515 161.405 ;
        RECT 21.980 161.110 24.515 161.250 ;
        RECT 27.070 161.250 27.390 161.310 ;
        RECT 28.910 161.250 29.230 161.310 ;
        RECT 27.070 161.110 29.230 161.250 ;
        RECT 21.980 161.065 22.270 161.110 ;
        RECT 27.070 161.050 27.390 161.110 ;
        RECT 28.910 161.050 29.230 161.110 ;
        RECT 25.245 160.910 25.535 160.955 ;
        RECT 25.690 160.910 26.010 160.970 ;
        RECT 25.245 160.770 26.010 160.910 ;
        RECT 25.245 160.725 25.535 160.770 ;
        RECT 25.690 160.710 26.010 160.770 ;
        RECT 21.980 160.570 22.270 160.615 ;
        RECT 24.760 160.570 25.050 160.615 ;
        RECT 26.620 160.570 26.910 160.615 ;
        RECT 21.980 160.430 26.910 160.570 ;
        RECT 21.980 160.385 22.270 160.430 ;
        RECT 24.760 160.385 25.050 160.430 ;
        RECT 26.620 160.385 26.910 160.430 ;
        RECT 29.460 160.570 29.600 161.405 ;
        RECT 31.210 161.390 31.530 161.450 ;
        RECT 34.905 161.405 35.195 161.450 ;
        RECT 35.365 161.405 35.655 161.635 ;
        RECT 36.270 161.590 36.590 161.650 ;
        RECT 45.945 161.590 46.235 161.635 ;
        RECT 49.700 161.590 49.840 161.730 ;
        RECT 36.270 161.450 46.235 161.590 ;
        RECT 33.970 161.250 34.290 161.310 ;
        RECT 35.440 161.250 35.580 161.405 ;
        RECT 36.270 161.390 36.590 161.450 ;
        RECT 45.945 161.405 46.235 161.450 ;
        RECT 49.240 161.450 49.840 161.590 ;
        RECT 43.185 161.250 43.475 161.295 ;
        RECT 48.705 161.250 48.995 161.295 ;
        RECT 33.970 161.110 35.580 161.250 ;
        RECT 40.040 161.110 41.100 161.250 ;
        RECT 33.970 161.050 34.290 161.110 ;
        RECT 30.750 160.910 31.070 160.970 ;
        RECT 36.285 160.910 36.575 160.955 ;
        RECT 40.040 160.910 40.180 161.110 ;
        RECT 30.750 160.770 40.180 160.910 ;
        RECT 30.750 160.710 31.070 160.770 ;
        RECT 36.285 160.725 36.575 160.770 ;
        RECT 40.425 160.725 40.715 160.955 ;
        RECT 40.960 160.910 41.100 161.110 ;
        RECT 43.185 161.110 48.995 161.250 ;
        RECT 43.185 161.065 43.475 161.110 ;
        RECT 48.705 161.065 48.995 161.110 ;
        RECT 49.240 160.970 49.380 161.450 ;
        RECT 49.610 161.250 49.930 161.310 ;
        RECT 51.005 161.250 51.295 161.295 ;
        RECT 54.685 161.250 54.975 161.295 ;
        RECT 49.610 161.110 54.975 161.250 ;
        RECT 57.060 161.250 57.200 161.745 ;
        RECT 62.490 161.730 62.810 161.790 ;
        RECT 82.730 161.930 83.050 161.990 ;
        RECT 89.875 161.930 90.165 161.975 ;
        RECT 94.690 161.930 95.010 161.990 ;
        RECT 82.730 161.790 84.340 161.930 ;
        RECT 82.730 161.730 83.050 161.790 ;
        RECT 84.200 161.635 84.340 161.790 ;
        RECT 87.880 161.790 95.010 161.930 ;
        RECT 84.125 161.590 84.415 161.635 ;
        RECT 87.880 161.590 88.020 161.790 ;
        RECT 89.875 161.745 90.165 161.790 ;
        RECT 94.690 161.730 95.010 161.790 ;
        RECT 105.745 161.930 106.035 161.975 ;
        RECT 106.190 161.930 106.510 161.990 ;
        RECT 105.745 161.790 106.510 161.930 ;
        RECT 105.745 161.745 106.035 161.790 ;
        RECT 106.190 161.730 106.510 161.790 ;
        RECT 109.870 161.930 110.190 161.990 ;
        RECT 111.725 161.930 112.015 161.975 ;
        RECT 109.870 161.790 112.015 161.930 ;
        RECT 109.870 161.730 110.190 161.790 ;
        RECT 111.725 161.745 112.015 161.790 ;
        RECT 114.025 161.745 114.315 161.975 ;
        RECT 116.310 161.930 116.630 161.990 ;
        RECT 116.785 161.930 117.075 161.975 ;
        RECT 117.230 161.930 117.550 161.990 ;
        RECT 116.310 161.790 117.550 161.930 ;
        RECT 68.100 161.450 70.540 161.590 ;
        RECT 59.745 161.250 60.035 161.295 ;
        RECT 57.060 161.110 60.035 161.250 ;
        RECT 49.610 161.050 49.930 161.110 ;
        RECT 51.005 161.065 51.295 161.110 ;
        RECT 54.685 161.065 54.975 161.110 ;
        RECT 59.745 161.065 60.035 161.110 ;
        RECT 66.185 161.250 66.475 161.295 ;
        RECT 66.630 161.250 66.950 161.310 ;
        RECT 68.100 161.295 68.240 161.450 ;
        RECT 70.400 161.295 70.540 161.450 ;
        RECT 84.125 161.450 88.020 161.590 ;
        RECT 91.880 161.590 92.170 161.635 ;
        RECT 94.230 161.590 94.550 161.650 ;
        RECT 95.140 161.590 95.430 161.635 ;
        RECT 91.880 161.450 95.430 161.590 ;
        RECT 84.125 161.405 84.415 161.450 ;
        RECT 91.880 161.405 92.170 161.450 ;
        RECT 94.230 161.390 94.550 161.450 ;
        RECT 95.140 161.405 95.430 161.450 ;
        RECT 96.060 161.590 96.350 161.635 ;
        RECT 97.920 161.590 98.210 161.635 ;
        RECT 96.060 161.450 98.210 161.590 ;
        RECT 114.100 161.590 114.240 161.745 ;
        RECT 116.310 161.730 116.630 161.790 ;
        RECT 116.785 161.745 117.075 161.790 ;
        RECT 117.230 161.730 117.550 161.790 ;
        RECT 119.530 161.730 119.850 161.990 ;
        RECT 121.370 161.930 121.690 161.990 ;
        RECT 121.845 161.930 122.135 161.975 ;
        RECT 121.370 161.790 122.135 161.930 ;
        RECT 121.370 161.730 121.690 161.790 ;
        RECT 121.845 161.745 122.135 161.790 ;
        RECT 123.670 161.590 123.990 161.650 ;
        RECT 114.100 161.450 123.990 161.590 ;
        RECT 96.060 161.405 96.350 161.450 ;
        RECT 97.920 161.405 98.210 161.450 ;
        RECT 66.185 161.110 67.780 161.250 ;
        RECT 66.185 161.065 66.475 161.110 ;
        RECT 66.630 161.050 66.950 161.110 ;
        RECT 46.865 160.910 47.155 160.955 ;
        RECT 40.960 160.770 47.155 160.910 ;
        RECT 46.865 160.725 47.155 160.770 ;
        RECT 49.150 160.910 49.470 160.970 ;
        RECT 51.465 160.910 51.755 160.955 ;
        RECT 49.150 160.770 51.755 160.910 ;
        RECT 37.650 160.570 37.970 160.630 ;
        RECT 29.460 160.430 37.970 160.570 ;
        RECT 40.500 160.570 40.640 160.725 ;
        RECT 43.645 160.570 43.935 160.615 ;
        RECT 40.500 160.430 43.935 160.570 ;
        RECT 46.940 160.570 47.080 160.725 ;
        RECT 49.150 160.710 49.470 160.770 ;
        RECT 51.465 160.725 51.755 160.770 ;
        RECT 52.385 160.910 52.675 160.955 ;
        RECT 54.225 160.910 54.515 160.955 ;
        RECT 67.090 160.910 67.410 160.970 ;
        RECT 52.385 160.770 67.410 160.910 ;
        RECT 67.640 160.910 67.780 161.110 ;
        RECT 68.025 161.065 68.315 161.295 ;
        RECT 68.485 161.065 68.775 161.295 ;
        RECT 70.325 161.250 70.615 161.295 ;
        RECT 71.230 161.250 71.550 161.310 ;
        RECT 70.325 161.110 71.550 161.250 ;
        RECT 70.325 161.065 70.615 161.110 ;
        RECT 68.560 160.910 68.700 161.065 ;
        RECT 71.230 161.050 71.550 161.110 ;
        RECT 81.825 161.250 82.115 161.295 ;
        RECT 86.425 161.250 86.715 161.295 ;
        RECT 81.825 161.110 85.720 161.250 ;
        RECT 81.825 161.065 82.115 161.110 ;
        RECT 67.640 160.770 68.700 160.910 ;
        RECT 79.970 160.910 80.290 160.970 ;
        RECT 82.745 160.910 83.035 160.955 ;
        RECT 79.970 160.770 83.035 160.910 ;
        RECT 52.385 160.725 52.675 160.770 ;
        RECT 54.225 160.725 54.515 160.770 ;
        RECT 52.460 160.570 52.600 160.725 ;
        RECT 67.090 160.710 67.410 160.770 ;
        RECT 79.970 160.710 80.290 160.770 ;
        RECT 82.745 160.725 83.035 160.770 ;
        RECT 83.665 160.725 83.955 160.955 ;
        RECT 46.940 160.430 52.600 160.570 ;
        RECT 53.290 160.570 53.610 160.630 ;
        RECT 65.265 160.570 65.555 160.615 ;
        RECT 70.770 160.570 71.090 160.630 ;
        RECT 53.290 160.430 71.090 160.570 ;
        RECT 18.115 160.230 18.405 160.275 ;
        RECT 21.550 160.230 21.870 160.290 ;
        RECT 29.460 160.230 29.600 160.430 ;
        RECT 37.650 160.370 37.970 160.430 ;
        RECT 43.645 160.385 43.935 160.430 ;
        RECT 53.290 160.370 53.610 160.430 ;
        RECT 65.265 160.385 65.555 160.430 ;
        RECT 70.770 160.370 71.090 160.430 ;
        RECT 80.890 160.570 81.210 160.630 ;
        RECT 83.740 160.570 83.880 160.725 ;
        RECT 80.890 160.430 83.880 160.570 ;
        RECT 80.890 160.370 81.210 160.430 ;
        RECT 18.115 160.090 29.600 160.230 ;
        RECT 33.970 160.230 34.290 160.290 ;
        RECT 34.890 160.230 35.210 160.290 ;
        RECT 33.970 160.090 35.210 160.230 ;
        RECT 18.115 160.045 18.405 160.090 ;
        RECT 21.550 160.030 21.870 160.090 ;
        RECT 33.970 160.030 34.290 160.090 ;
        RECT 34.890 160.030 35.210 160.090 ;
        RECT 67.090 160.030 67.410 160.290 ;
        RECT 69.405 160.230 69.695 160.275 ;
        RECT 69.850 160.230 70.170 160.290 ;
        RECT 69.405 160.090 70.170 160.230 ;
        RECT 69.405 160.045 69.695 160.090 ;
        RECT 69.850 160.030 70.170 160.090 ;
        RECT 71.245 160.230 71.535 160.275 ;
        RECT 73.990 160.230 74.310 160.290 ;
        RECT 71.245 160.090 74.310 160.230 ;
        RECT 71.245 160.045 71.535 160.090 ;
        RECT 73.990 160.030 74.310 160.090 ;
        RECT 81.365 160.230 81.655 160.275 ;
        RECT 83.190 160.230 83.510 160.290 ;
        RECT 81.365 160.090 83.510 160.230 ;
        RECT 85.580 160.230 85.720 161.110 ;
        RECT 86.040 161.110 86.715 161.250 ;
        RECT 86.040 160.615 86.180 161.110 ;
        RECT 86.425 161.065 86.715 161.110 ;
        RECT 93.740 161.250 94.030 161.295 ;
        RECT 96.060 161.250 96.275 161.405 ;
        RECT 123.670 161.390 123.990 161.450 ;
        RECT 93.740 161.110 96.275 161.250 ;
        RECT 97.450 161.250 97.770 161.310 ;
        RECT 98.845 161.250 99.135 161.295 ;
        RECT 102.065 161.250 102.355 161.295 ;
        RECT 97.450 161.110 102.355 161.250 ;
        RECT 93.740 161.065 94.030 161.110 ;
        RECT 97.450 161.050 97.770 161.110 ;
        RECT 98.845 161.065 99.135 161.110 ;
        RECT 102.065 161.065 102.355 161.110 ;
        RECT 96.990 160.710 97.310 160.970 ;
        RECT 102.140 160.910 102.280 161.065 ;
        RECT 102.510 161.050 102.830 161.310 ;
        RECT 107.125 161.250 107.415 161.295 ;
        RECT 110.330 161.250 110.650 161.310 ;
        RECT 107.125 161.110 110.650 161.250 ;
        RECT 107.125 161.065 107.415 161.110 ;
        RECT 110.330 161.050 110.650 161.110 ;
        RECT 112.185 161.250 112.475 161.295 ;
        RECT 114.010 161.250 114.330 161.310 ;
        RECT 116.325 161.250 116.615 161.295 ;
        RECT 112.185 161.110 116.615 161.250 ;
        RECT 112.185 161.065 112.475 161.110 ;
        RECT 114.010 161.050 114.330 161.110 ;
        RECT 116.325 161.065 116.615 161.110 ;
        RECT 119.070 161.050 119.390 161.310 ;
        RECT 120.910 161.050 121.230 161.310 ;
        RECT 105.730 160.910 106.050 160.970 ;
        RECT 102.140 160.770 106.050 160.910 ;
        RECT 105.730 160.710 106.050 160.770 ;
        RECT 85.965 160.385 86.255 160.615 ;
        RECT 88.710 160.570 89.030 160.630 ;
        RECT 86.500 160.430 89.030 160.570 ;
        RECT 86.500 160.230 86.640 160.430 ;
        RECT 88.710 160.370 89.030 160.430 ;
        RECT 93.740 160.570 94.030 160.615 ;
        RECT 96.520 160.570 96.810 160.615 ;
        RECT 98.380 160.570 98.670 160.615 ;
        RECT 93.740 160.430 98.670 160.570 ;
        RECT 93.740 160.385 94.030 160.430 ;
        RECT 96.520 160.385 96.810 160.430 ;
        RECT 98.380 160.385 98.670 160.430 ;
        RECT 85.580 160.090 86.640 160.230 ;
        RECT 87.345 160.230 87.635 160.275 ;
        RECT 88.250 160.230 88.570 160.290 ;
        RECT 87.345 160.090 88.570 160.230 ;
        RECT 110.420 160.230 110.560 161.050 ;
        RECT 111.265 160.910 111.555 160.955 ;
        RECT 112.630 160.910 112.950 160.970 ;
        RECT 115.405 160.910 115.695 160.955 ;
        RECT 111.265 160.770 115.695 160.910 ;
        RECT 111.265 160.725 111.555 160.770 ;
        RECT 112.630 160.710 112.950 160.770 ;
        RECT 115.405 160.725 115.695 160.770 ;
        RECT 110.790 160.230 111.110 160.290 ;
        RECT 110.420 160.090 111.110 160.230 ;
        RECT 81.365 160.045 81.655 160.090 ;
        RECT 83.190 160.030 83.510 160.090 ;
        RECT 87.345 160.045 87.635 160.090 ;
        RECT 88.250 160.030 88.570 160.090 ;
        RECT 110.790 160.030 111.110 160.090 ;
        RECT 116.770 160.230 117.090 160.290 ;
        RECT 118.625 160.230 118.915 160.275 ;
        RECT 116.770 160.090 118.915 160.230 ;
        RECT 116.770 160.030 117.090 160.090 ;
        RECT 118.625 160.045 118.915 160.090 ;
        RECT 14.580 159.410 127.740 159.890 ;
        RECT 17.885 159.210 18.175 159.255 ;
        RECT 18.790 159.210 19.110 159.270 ;
        RECT 17.885 159.070 19.110 159.210 ;
        RECT 17.885 159.025 18.175 159.070 ;
        RECT 18.790 159.010 19.110 159.070 ;
        RECT 25.690 159.010 26.010 159.270 ;
        RECT 31.210 159.010 31.530 159.270 ;
        RECT 49.610 159.010 49.930 159.270 ;
        RECT 50.530 159.210 50.850 159.270 ;
        RECT 52.830 159.210 53.150 159.270 ;
        RECT 50.530 159.070 53.150 159.210 ;
        RECT 50.530 159.010 50.850 159.070 ;
        RECT 52.830 159.010 53.150 159.070 ;
        RECT 71.245 159.210 71.535 159.255 ;
        RECT 71.690 159.210 72.010 159.270 ;
        RECT 71.245 159.070 72.010 159.210 ;
        RECT 71.245 159.025 71.535 159.070 ;
        RECT 71.690 159.010 72.010 159.070 ;
        RECT 79.970 159.010 80.290 159.270 ;
        RECT 80.890 159.255 81.210 159.270 ;
        RECT 80.890 159.025 81.425 159.255 ;
        RECT 93.325 159.210 93.615 159.255 ;
        RECT 94.230 159.210 94.550 159.270 ;
        RECT 93.325 159.070 94.550 159.210 ;
        RECT 93.325 159.025 93.615 159.070 ;
        RECT 80.890 159.010 81.210 159.025 ;
        RECT 94.230 159.010 94.550 159.070 ;
        RECT 96.990 159.210 97.310 159.270 ;
        RECT 97.465 159.210 97.755 159.255 ;
        RECT 96.990 159.070 97.755 159.210 ;
        RECT 96.990 159.010 97.310 159.070 ;
        RECT 97.465 159.025 97.755 159.070 ;
        RECT 100.210 159.010 100.530 159.270 ;
        RECT 104.365 159.210 104.655 159.255 ;
        RECT 104.810 159.210 105.130 159.270 ;
        RECT 112.170 159.210 112.490 159.270 ;
        RECT 104.365 159.070 105.130 159.210 ;
        RECT 104.365 159.025 104.655 159.070 ;
        RECT 104.810 159.010 105.130 159.070 ;
        RECT 110.420 159.070 112.490 159.210 ;
        RECT 30.750 158.870 31.070 158.930 ;
        RECT 21.180 158.730 31.070 158.870 ;
        RECT 21.180 158.590 21.320 158.730 ;
        RECT 30.750 158.670 31.070 158.730 ;
        RECT 42.570 158.730 53.980 158.870 ;
        RECT 21.090 158.330 21.410 158.590 ;
        RECT 21.550 158.330 21.870 158.590 ;
        RECT 29.830 158.530 30.150 158.590 ;
        RECT 42.570 158.530 42.710 158.730 ;
        RECT 22.790 158.390 30.150 158.530 ;
        RECT 18.345 158.190 18.635 158.235 ;
        RECT 18.805 158.190 19.095 158.235 ;
        RECT 22.790 158.190 22.930 158.390 ;
        RECT 29.830 158.330 30.150 158.390 ;
        RECT 39.120 158.390 42.710 158.530 ;
        RECT 24.785 158.190 25.075 158.235 ;
        RECT 18.345 158.050 22.930 158.190 ;
        RECT 23.940 158.050 25.075 158.190 ;
        RECT 18.345 158.005 18.635 158.050 ;
        RECT 18.805 158.005 19.095 158.050 ;
        RECT 19.250 157.310 19.570 157.570 ;
        RECT 22.010 157.310 22.330 157.570 ;
        RECT 23.940 157.555 24.080 158.050 ;
        RECT 24.785 158.005 25.075 158.050 ;
        RECT 28.465 158.005 28.755 158.235 ;
        RECT 32.130 158.190 32.450 158.250 ;
        RECT 35.810 158.190 36.130 158.250 ;
        RECT 39.120 158.235 39.260 158.390 ;
        RECT 32.130 158.050 36.130 158.190 ;
        RECT 28.540 157.850 28.680 158.005 ;
        RECT 32.130 157.990 32.450 158.050 ;
        RECT 35.810 157.990 36.130 158.050 ;
        RECT 39.045 158.005 39.335 158.235 ;
        RECT 39.965 158.005 40.255 158.235 ;
        RECT 40.425 158.005 40.715 158.235 ;
        RECT 40.885 158.190 41.175 158.235 ;
        RECT 41.790 158.190 42.110 158.250 ;
        RECT 40.885 158.050 42.110 158.190 ;
        RECT 42.570 158.235 42.710 158.390 ;
        RECT 46.865 158.530 47.155 158.575 ;
        RECT 50.530 158.530 50.850 158.590 ;
        RECT 53.840 158.530 53.980 158.730 ;
        RECT 69.405 158.685 69.695 158.915 ;
        RECT 70.770 158.870 71.090 158.930 ;
        RECT 85.000 158.870 85.290 158.915 ;
        RECT 87.780 158.870 88.070 158.915 ;
        RECT 89.640 158.870 89.930 158.915 ;
        RECT 70.770 158.730 78.360 158.870 ;
        RECT 69.480 158.530 69.620 158.685 ;
        RECT 70.770 158.670 71.090 158.730 ;
        RECT 46.865 158.390 50.850 158.530 ;
        RECT 46.865 158.345 47.155 158.390 ;
        RECT 50.530 158.330 50.850 158.390 ;
        RECT 52.000 158.390 53.520 158.530 ;
        RECT 42.570 158.050 42.955 158.235 ;
        RECT 40.885 158.005 41.175 158.050 ;
        RECT 36.270 157.850 36.590 157.910 ;
        RECT 40.040 157.850 40.180 158.005 ;
        RECT 28.540 157.710 40.180 157.850 ;
        RECT 40.500 157.850 40.640 158.005 ;
        RECT 41.790 157.990 42.110 158.050 ;
        RECT 42.665 158.005 42.955 158.050 ;
        RECT 43.170 158.190 43.490 158.250 ;
        RECT 43.645 158.190 43.935 158.235 ;
        RECT 43.170 158.050 43.935 158.190 ;
        RECT 43.170 157.990 43.490 158.050 ;
        RECT 43.645 158.005 43.935 158.050 ;
        RECT 44.105 158.005 44.395 158.235 ;
        RECT 44.565 158.190 44.855 158.235 ;
        RECT 45.010 158.190 45.330 158.250 ;
        RECT 52.000 158.235 52.140 158.390 ;
        RECT 51.925 158.190 52.215 158.235 ;
        RECT 44.565 158.050 52.215 158.190 ;
        RECT 44.565 158.005 44.855 158.050 ;
        RECT 44.180 157.850 44.320 158.005 ;
        RECT 45.010 157.990 45.330 158.050 ;
        RECT 51.925 158.005 52.215 158.050 ;
        RECT 52.385 158.005 52.675 158.235 ;
        RECT 52.460 157.850 52.600 158.005 ;
        RECT 52.830 157.990 53.150 158.250 ;
        RECT 40.500 157.710 52.600 157.850 ;
        RECT 53.380 157.850 53.520 158.390 ;
        RECT 53.840 158.390 72.380 158.530 ;
        RECT 53.840 158.250 53.980 158.390 ;
        RECT 53.750 157.990 54.070 158.250 ;
        RECT 56.970 158.190 57.290 158.250 ;
        RECT 61.125 158.190 61.415 158.235 ;
        RECT 62.505 158.190 62.795 158.235 ;
        RECT 56.970 158.050 62.795 158.190 ;
        RECT 56.970 157.990 57.290 158.050 ;
        RECT 61.125 158.005 61.415 158.050 ;
        RECT 62.505 158.005 62.795 158.050 ;
        RECT 62.950 158.190 63.270 158.250 ;
        RECT 63.885 158.190 64.175 158.235 ;
        RECT 62.950 158.050 64.175 158.190 ;
        RECT 62.950 157.990 63.270 158.050 ;
        RECT 63.885 158.005 64.175 158.050 ;
        RECT 68.485 158.190 68.775 158.235 ;
        RECT 69.390 158.190 69.710 158.250 ;
        RECT 70.310 158.190 70.630 158.250 ;
        RECT 72.240 158.235 72.380 158.390 ;
        RECT 68.485 158.050 70.630 158.190 ;
        RECT 68.485 158.005 68.775 158.050 ;
        RECT 69.390 157.990 69.710 158.050 ;
        RECT 70.310 157.990 70.630 158.050 ;
        RECT 72.165 158.005 72.455 158.235 ;
        RECT 72.240 157.850 72.380 158.005 ;
        RECT 73.070 157.990 73.390 158.250 ;
        RECT 73.620 158.235 73.760 158.730 ;
        RECT 76.290 158.530 76.610 158.590 ;
        RECT 76.290 158.390 77.900 158.530 ;
        RECT 76.290 158.330 76.610 158.390 ;
        RECT 73.545 158.005 73.835 158.235 ;
        RECT 73.990 157.990 74.310 158.250 ;
        RECT 77.760 158.235 77.900 158.390 ;
        RECT 78.220 158.235 78.360 158.730 ;
        RECT 85.000 158.730 89.930 158.870 ;
        RECT 85.000 158.685 85.290 158.730 ;
        RECT 87.780 158.685 88.070 158.730 ;
        RECT 89.640 158.685 89.930 158.730 ;
        RECT 106.665 158.870 106.955 158.915 ;
        RECT 109.410 158.870 109.730 158.930 ;
        RECT 106.665 158.730 109.730 158.870 ;
        RECT 106.665 158.685 106.955 158.730 ;
        RECT 109.410 158.670 109.730 158.730 ;
        RECT 88.250 158.330 88.570 158.590 ;
        RECT 88.710 158.530 89.030 158.590 ;
        RECT 88.710 158.390 93.080 158.530 ;
        RECT 88.710 158.330 89.030 158.390 ;
        RECT 76.765 158.190 77.055 158.235 ;
        RECT 76.380 158.050 77.055 158.190 ;
        RECT 76.380 157.910 76.520 158.050 ;
        RECT 76.765 158.005 77.055 158.050 ;
        RECT 77.685 158.005 77.975 158.235 ;
        RECT 78.145 158.005 78.435 158.235 ;
        RECT 78.605 158.190 78.895 158.235 ;
        RECT 79.050 158.190 79.370 158.250 ;
        RECT 81.810 158.190 82.130 158.250 ;
        RECT 78.605 158.050 82.130 158.190 ;
        RECT 78.605 158.005 78.895 158.050 ;
        RECT 76.290 157.850 76.610 157.910 ;
        RECT 53.380 157.710 61.340 157.850 ;
        RECT 72.240 157.710 76.610 157.850 ;
        RECT 78.220 157.850 78.360 158.005 ;
        RECT 79.050 157.990 79.370 158.050 ;
        RECT 81.810 157.990 82.130 158.050 ;
        RECT 85.000 158.190 85.290 158.235 ;
        RECT 90.105 158.190 90.395 158.235 ;
        RECT 91.010 158.190 91.330 158.250 ;
        RECT 92.940 158.235 93.080 158.390 ;
        RECT 85.000 158.050 87.535 158.190 ;
        RECT 85.000 158.005 85.290 158.050 ;
        RECT 82.270 157.850 82.590 157.910 ;
        RECT 83.190 157.895 83.510 157.910 ;
        RECT 87.320 157.895 87.535 158.050 ;
        RECT 90.105 158.050 91.330 158.190 ;
        RECT 90.105 158.005 90.395 158.050 ;
        RECT 91.010 157.990 91.330 158.050 ;
        RECT 92.865 158.005 93.155 158.235 ;
        RECT 78.220 157.710 82.590 157.850 ;
        RECT 36.270 157.650 36.590 157.710 ;
        RECT 43.260 157.570 43.400 157.710 ;
        RECT 23.865 157.325 24.155 157.555 ;
        RECT 34.890 157.310 35.210 157.570 ;
        RECT 42.250 157.310 42.570 157.570 ;
        RECT 43.170 157.310 43.490 157.570 ;
        RECT 45.930 157.310 46.250 157.570 ;
        RECT 50.070 157.510 50.390 157.570 ;
        RECT 50.545 157.510 50.835 157.555 ;
        RECT 50.070 157.370 50.835 157.510 ;
        RECT 52.460 157.510 52.600 157.710 ;
        RECT 53.290 157.510 53.610 157.570 ;
        RECT 52.460 157.370 53.610 157.510 ;
        RECT 50.070 157.310 50.390 157.370 ;
        RECT 50.545 157.325 50.835 157.370 ;
        RECT 53.290 157.310 53.610 157.370 ;
        RECT 58.810 157.510 59.130 157.570 ;
        RECT 60.665 157.510 60.955 157.555 ;
        RECT 58.810 157.370 60.955 157.510 ;
        RECT 61.200 157.510 61.340 157.710 ;
        RECT 76.290 157.650 76.610 157.710 ;
        RECT 82.270 157.650 82.590 157.710 ;
        RECT 83.140 157.850 83.510 157.895 ;
        RECT 86.400 157.850 86.690 157.895 ;
        RECT 83.140 157.710 86.690 157.850 ;
        RECT 83.140 157.665 83.510 157.710 ;
        RECT 86.400 157.665 86.690 157.710 ;
        RECT 87.320 157.850 87.610 157.895 ;
        RECT 89.180 157.850 89.470 157.895 ;
        RECT 87.320 157.710 89.470 157.850 ;
        RECT 92.940 157.850 93.080 158.005 ;
        RECT 96.530 157.990 96.850 158.250 ;
        RECT 99.765 158.005 100.055 158.235 ;
        RECT 95.150 157.850 95.470 157.910 ;
        RECT 99.840 157.850 99.980 158.005 ;
        RECT 105.270 157.990 105.590 158.250 ;
        RECT 105.745 158.190 106.035 158.235 ;
        RECT 108.950 158.190 109.270 158.250 ;
        RECT 105.745 158.050 109.270 158.190 ;
        RECT 105.745 158.005 106.035 158.050 ;
        RECT 108.950 157.990 109.270 158.050 ;
        RECT 109.410 157.990 109.730 158.250 ;
        RECT 109.870 157.990 110.190 158.250 ;
        RECT 110.420 158.235 110.560 159.070 ;
        RECT 112.170 159.010 112.490 159.070 ;
        RECT 119.545 159.210 119.835 159.255 ;
        RECT 120.910 159.210 121.230 159.270 ;
        RECT 119.545 159.070 121.230 159.210 ;
        RECT 119.545 159.025 119.835 159.070 ;
        RECT 120.910 159.010 121.230 159.070 ;
        RECT 116.770 158.330 117.090 158.590 ;
        RECT 110.345 158.005 110.635 158.235 ;
        RECT 111.265 158.190 111.555 158.235 ;
        RECT 111.710 158.190 112.030 158.250 ;
        RECT 111.265 158.050 112.030 158.190 ;
        RECT 111.265 158.005 111.555 158.050 ;
        RECT 111.710 157.990 112.030 158.050 ;
        RECT 112.170 157.850 112.490 157.910 ;
        RECT 92.940 157.710 112.490 157.850 ;
        RECT 87.320 157.665 87.610 157.710 ;
        RECT 89.180 157.665 89.470 157.710 ;
        RECT 83.190 157.650 83.510 157.665 ;
        RECT 95.150 157.650 95.470 157.710 ;
        RECT 112.170 157.650 112.490 157.710 ;
        RECT 73.990 157.510 74.310 157.570 ;
        RECT 61.200 157.370 74.310 157.510 ;
        RECT 58.810 157.310 59.130 157.370 ;
        RECT 60.665 157.325 60.955 157.370 ;
        RECT 73.990 157.310 74.310 157.370 ;
        RECT 75.385 157.510 75.675 157.555 ;
        RECT 75.830 157.510 76.150 157.570 ;
        RECT 75.385 157.370 76.150 157.510 ;
        RECT 75.385 157.325 75.675 157.370 ;
        RECT 75.830 157.310 76.150 157.370 ;
        RECT 108.045 157.510 108.335 157.555 ;
        RECT 108.950 157.510 109.270 157.570 ;
        RECT 108.045 157.370 109.270 157.510 ;
        RECT 108.045 157.325 108.335 157.370 ;
        RECT 108.950 157.310 109.270 157.370 ;
        RECT 14.580 156.690 127.740 157.170 ;
        RECT 17.195 156.490 17.485 156.535 ;
        RECT 22.010 156.490 22.330 156.550 ;
        RECT 33.510 156.490 33.830 156.550 ;
        RECT 34.445 156.490 34.735 156.535 ;
        RECT 17.195 156.350 32.820 156.490 ;
        RECT 17.195 156.305 17.485 156.350 ;
        RECT 22.010 156.290 22.330 156.350 ;
        RECT 19.250 156.195 19.570 156.210 ;
        RECT 19.200 156.150 19.570 156.195 ;
        RECT 22.460 156.150 22.750 156.195 ;
        RECT 19.200 156.010 22.750 156.150 ;
        RECT 19.200 155.965 19.570 156.010 ;
        RECT 22.460 155.965 22.750 156.010 ;
        RECT 23.380 156.150 23.670 156.195 ;
        RECT 25.240 156.150 25.530 156.195 ;
        RECT 23.380 156.010 25.530 156.150 ;
        RECT 32.680 156.150 32.820 156.350 ;
        RECT 33.510 156.350 34.735 156.490 ;
        RECT 33.510 156.290 33.830 156.350 ;
        RECT 34.445 156.305 34.735 156.350 ;
        RECT 34.890 156.290 35.210 156.550 ;
        RECT 41.790 156.490 42.110 156.550 ;
        RECT 45.010 156.490 45.330 156.550 ;
        RECT 40.500 156.350 45.330 156.490 ;
        RECT 32.680 156.010 34.660 156.150 ;
        RECT 23.380 155.965 23.670 156.010 ;
        RECT 25.240 155.965 25.530 156.010 ;
        RECT 19.250 155.950 19.570 155.965 ;
        RECT 21.060 155.810 21.350 155.855 ;
        RECT 23.380 155.810 23.595 155.965 ;
        RECT 21.060 155.670 23.595 155.810 ;
        RECT 26.165 155.810 26.455 155.855 ;
        RECT 27.070 155.810 27.390 155.870 ;
        RECT 26.165 155.670 27.390 155.810 ;
        RECT 21.060 155.625 21.350 155.670 ;
        RECT 26.165 155.625 26.455 155.670 ;
        RECT 27.070 155.610 27.390 155.670 ;
        RECT 27.530 155.610 27.850 155.870 ;
        RECT 31.210 155.810 31.530 155.870 ;
        RECT 33.510 155.810 33.830 155.870 ;
        RECT 31.210 155.670 33.830 155.810 ;
        RECT 31.210 155.610 31.530 155.670 ;
        RECT 33.510 155.610 33.830 155.670 ;
        RECT 24.325 155.470 24.615 155.515 ;
        RECT 30.750 155.470 31.070 155.530 ;
        RECT 33.970 155.470 34.290 155.530 ;
        RECT 24.325 155.330 26.840 155.470 ;
        RECT 24.325 155.285 24.615 155.330 ;
        RECT 26.700 155.175 26.840 155.330 ;
        RECT 30.750 155.330 34.290 155.470 ;
        RECT 34.520 155.470 34.660 156.010 ;
        RECT 40.500 155.810 40.640 156.350 ;
        RECT 41.790 156.290 42.110 156.350 ;
        RECT 45.010 156.290 45.330 156.350 ;
        RECT 49.150 156.490 49.470 156.550 ;
        RECT 50.530 156.490 50.850 156.550 ;
        RECT 67.090 156.490 67.410 156.550 ;
        RECT 102.510 156.490 102.830 156.550 ;
        RECT 108.490 156.490 108.810 156.550 ;
        RECT 111.710 156.490 112.030 156.550 ;
        RECT 49.150 156.350 49.840 156.490 ;
        RECT 49.150 156.290 49.470 156.350 ;
        RECT 40.870 156.150 41.190 156.210 ;
        RECT 45.100 156.150 45.240 156.290 ;
        RECT 40.870 156.010 43.400 156.150 ;
        RECT 40.870 155.950 41.190 156.010 ;
        RECT 41.345 155.810 41.635 155.855 ;
        RECT 40.500 155.670 41.635 155.810 ;
        RECT 41.345 155.625 41.635 155.670 ;
        RECT 41.790 155.610 42.110 155.870 ;
        RECT 43.260 155.855 43.400 156.010 ;
        RECT 45.100 156.010 48.920 156.150 ;
        RECT 45.100 155.855 45.240 156.010 ;
        RECT 42.265 155.625 42.555 155.855 ;
        RECT 43.185 155.625 43.475 155.855 ;
        RECT 45.025 155.625 45.315 155.855 ;
        RECT 45.470 155.625 45.760 155.855 ;
        RECT 45.970 155.625 46.260 155.855 ;
        RECT 42.340 155.470 42.480 155.625 ;
        RECT 34.520 155.330 42.480 155.470 ;
        RECT 43.630 155.470 43.950 155.530 ;
        RECT 45.560 155.470 45.700 155.625 ;
        RECT 43.630 155.330 45.700 155.470 ;
        RECT 30.750 155.270 31.070 155.330 ;
        RECT 33.970 155.270 34.290 155.330 ;
        RECT 43.630 155.270 43.950 155.330 ;
        RECT 21.060 155.130 21.350 155.175 ;
        RECT 23.840 155.130 24.130 155.175 ;
        RECT 25.700 155.130 25.990 155.175 ;
        RECT 21.060 154.990 25.990 155.130 ;
        RECT 21.060 154.945 21.350 154.990 ;
        RECT 23.840 154.945 24.130 154.990 ;
        RECT 25.700 154.945 25.990 154.990 ;
        RECT 26.625 154.945 26.915 155.175 ;
        RECT 32.130 155.130 32.450 155.190 ;
        RECT 46.020 155.130 46.160 155.625 ;
        RECT 46.850 155.610 47.170 155.870 ;
        RECT 48.780 155.855 48.920 156.010 ;
        RECT 49.700 155.855 49.840 156.350 ;
        RECT 50.530 156.350 85.030 156.490 ;
        RECT 50.530 156.290 50.850 156.350 ;
        RECT 67.090 156.290 67.410 156.350 ;
        RECT 53.290 156.150 53.610 156.210 ;
        RECT 58.810 156.195 59.130 156.210 ;
        RECT 50.160 156.010 53.610 156.150 ;
        RECT 48.705 155.625 48.995 155.855 ;
        RECT 49.165 155.625 49.455 155.855 ;
        RECT 49.625 155.625 49.915 155.855 ;
        RECT 49.240 155.470 49.380 155.625 ;
        RECT 50.160 155.470 50.300 156.010 ;
        RECT 53.290 155.950 53.610 156.010 ;
        RECT 55.540 156.150 55.830 156.195 ;
        RECT 58.800 156.150 59.130 156.195 ;
        RECT 55.540 156.010 59.130 156.150 ;
        RECT 55.540 155.965 55.830 156.010 ;
        RECT 58.800 155.965 59.130 156.010 ;
        RECT 58.810 155.950 59.130 155.965 ;
        RECT 59.720 156.150 60.010 156.195 ;
        RECT 61.580 156.150 61.870 156.195 ;
        RECT 59.720 156.010 61.870 156.150 ;
        RECT 59.720 155.965 60.010 156.010 ;
        RECT 61.580 155.965 61.870 156.010 ;
        RECT 73.990 156.150 74.310 156.210 ;
        RECT 80.890 156.150 81.210 156.210 ;
        RECT 73.990 156.010 78.360 156.150 ;
        RECT 50.545 155.810 50.835 155.855 ;
        RECT 53.750 155.810 54.070 155.870 ;
        RECT 50.545 155.670 54.070 155.810 ;
        RECT 50.545 155.625 50.835 155.670 ;
        RECT 49.240 155.330 50.300 155.470 ;
        RECT 32.130 154.990 46.160 155.130 ;
        RECT 46.850 155.130 47.170 155.190 ;
        RECT 50.620 155.130 50.760 155.625 ;
        RECT 53.750 155.610 54.070 155.670 ;
        RECT 57.400 155.810 57.690 155.855 ;
        RECT 59.720 155.810 59.935 155.965 ;
        RECT 73.990 155.950 74.310 156.010 ;
        RECT 78.220 155.870 78.360 156.010 ;
        RECT 79.600 156.010 81.210 156.150 ;
        RECT 84.890 156.150 85.030 156.350 ;
        RECT 102.510 156.350 112.030 156.490 ;
        RECT 102.510 156.290 102.830 156.350 ;
        RECT 102.970 156.150 103.290 156.210 ;
        RECT 84.890 156.010 98.140 156.150 ;
        RECT 57.400 155.670 59.935 155.810 ;
        RECT 62.505 155.810 62.795 155.855 ;
        RECT 63.870 155.810 64.190 155.870 ;
        RECT 62.505 155.670 64.190 155.810 ;
        RECT 57.400 155.625 57.690 155.670 ;
        RECT 62.505 155.625 62.795 155.670 ;
        RECT 63.870 155.610 64.190 155.670 ;
        RECT 74.450 155.610 74.770 155.870 ;
        RECT 78.130 155.610 78.450 155.870 ;
        RECT 78.590 155.610 78.910 155.870 ;
        RECT 79.065 155.810 79.355 155.855 ;
        RECT 79.600 155.810 79.740 156.010 ;
        RECT 80.890 155.950 81.210 156.010 ;
        RECT 79.065 155.670 79.740 155.810 ;
        RECT 79.065 155.625 79.355 155.670 ;
        RECT 79.985 155.625 80.275 155.855 ;
        RECT 60.665 155.470 60.955 155.515 ;
        RECT 61.110 155.470 61.430 155.530 ;
        RECT 60.665 155.330 61.430 155.470 ;
        RECT 60.665 155.285 60.955 155.330 ;
        RECT 61.110 155.270 61.430 155.330 ;
        RECT 65.710 155.270 66.030 155.530 ;
        RECT 76.290 155.470 76.610 155.530 ;
        RECT 80.060 155.470 80.200 155.625 ;
        RECT 81.810 155.610 82.130 155.870 ;
        RECT 82.270 155.610 82.590 155.870 ;
        RECT 82.730 155.610 83.050 155.870 ;
        RECT 83.665 155.625 83.955 155.855 ;
        RECT 84.570 155.810 84.890 155.870 ;
        RECT 97.465 155.810 97.755 155.855 ;
        RECT 84.570 155.670 97.755 155.810 ;
        RECT 83.740 155.470 83.880 155.625 ;
        RECT 84.570 155.610 84.890 155.670 ;
        RECT 97.465 155.625 97.755 155.670 ;
        RECT 76.290 155.330 83.880 155.470 ;
        RECT 76.290 155.270 76.610 155.330 ;
        RECT 46.850 154.990 50.760 155.130 ;
        RECT 57.400 155.130 57.690 155.175 ;
        RECT 60.180 155.130 60.470 155.175 ;
        RECT 62.040 155.130 62.330 155.175 ;
        RECT 57.400 154.990 62.330 155.130 ;
        RECT 32.130 154.930 32.450 154.990 ;
        RECT 46.850 154.930 47.170 154.990 ;
        RECT 57.400 154.945 57.690 154.990 ;
        RECT 60.180 154.945 60.470 154.990 ;
        RECT 62.040 154.945 62.330 154.990 ;
        RECT 78.590 155.130 78.910 155.190 ;
        RECT 82.270 155.130 82.590 155.190 ;
        RECT 78.590 154.990 82.590 155.130 ;
        RECT 97.540 155.130 97.680 155.625 ;
        RECT 98.000 155.470 98.140 156.010 ;
        RECT 102.970 156.010 106.420 156.150 ;
        RECT 102.970 155.950 103.290 156.010 ;
        RECT 98.370 155.610 98.690 155.870 ;
        RECT 98.830 155.610 99.150 155.870 ;
        RECT 99.305 155.810 99.595 155.855 ;
        RECT 104.825 155.810 105.115 155.855 ;
        RECT 99.305 155.670 105.115 155.810 ;
        RECT 99.305 155.625 99.595 155.670 ;
        RECT 104.825 155.625 105.115 155.670 ;
        RECT 99.380 155.470 99.520 155.625 ;
        RECT 98.000 155.330 99.520 155.470 ;
        RECT 102.510 155.130 102.830 155.190 ;
        RECT 97.540 154.990 102.830 155.130 ;
        RECT 78.590 154.930 78.910 154.990 ;
        RECT 82.270 154.930 82.590 154.990 ;
        RECT 102.510 154.930 102.830 154.990 ;
        RECT 35.810 154.790 36.130 154.850 ;
        RECT 36.745 154.790 37.035 154.835 ;
        RECT 35.810 154.650 37.035 154.790 ;
        RECT 35.810 154.590 36.130 154.650 ;
        RECT 36.745 154.605 37.035 154.650 ;
        RECT 39.950 154.590 40.270 154.850 ;
        RECT 43.630 154.590 43.950 154.850 ;
        RECT 45.010 154.790 45.330 154.850 ;
        RECT 46.940 154.790 47.080 154.930 ;
        RECT 45.010 154.650 47.080 154.790 ;
        RECT 47.325 154.790 47.615 154.835 ;
        RECT 49.150 154.790 49.470 154.850 ;
        RECT 53.750 154.835 54.070 154.850 ;
        RECT 47.325 154.650 49.470 154.790 ;
        RECT 45.010 154.590 45.330 154.650 ;
        RECT 47.325 154.605 47.615 154.650 ;
        RECT 49.150 154.590 49.470 154.650 ;
        RECT 53.535 154.605 54.070 154.835 ;
        RECT 53.750 154.590 54.070 154.605 ;
        RECT 54.210 154.790 54.530 154.850 ;
        RECT 69.850 154.790 70.170 154.850 ;
        RECT 54.210 154.650 70.170 154.790 ;
        RECT 54.210 154.590 54.530 154.650 ;
        RECT 69.850 154.590 70.170 154.650 ;
        RECT 76.290 154.790 76.610 154.850 ;
        RECT 76.765 154.790 77.055 154.835 ;
        RECT 76.290 154.650 77.055 154.790 ;
        RECT 76.290 154.590 76.610 154.650 ;
        RECT 76.765 154.605 77.055 154.650 ;
        RECT 80.430 154.590 80.750 154.850 ;
        RECT 99.750 154.790 100.070 154.850 ;
        RECT 100.685 154.790 100.975 154.835 ;
        RECT 99.750 154.650 100.975 154.790 ;
        RECT 99.750 154.590 100.070 154.650 ;
        RECT 100.685 154.605 100.975 154.650 ;
        RECT 103.445 154.790 103.735 154.835 ;
        RECT 103.890 154.790 104.210 154.850 ;
        RECT 103.445 154.650 104.210 154.790 ;
        RECT 104.900 154.790 105.040 155.625 ;
        RECT 105.270 155.610 105.590 155.870 ;
        RECT 105.745 155.810 106.035 155.855 ;
        RECT 106.280 155.810 106.420 156.010 ;
        RECT 106.740 155.855 106.880 156.350 ;
        RECT 108.490 156.290 108.810 156.350 ;
        RECT 111.710 156.290 112.030 156.350 ;
        RECT 110.790 156.150 111.110 156.210 ;
        RECT 108.120 156.010 111.110 156.150 ;
        RECT 108.120 155.855 108.260 156.010 ;
        RECT 110.790 155.950 111.110 156.010 ;
        RECT 105.745 155.670 106.420 155.810 ;
        RECT 106.665 155.810 106.955 155.855 ;
        RECT 107.125 155.810 107.415 155.855 ;
        RECT 106.665 155.670 107.415 155.810 ;
        RECT 105.745 155.625 106.035 155.670 ;
        RECT 106.665 155.625 106.955 155.670 ;
        RECT 107.125 155.625 107.415 155.670 ;
        RECT 108.045 155.625 108.335 155.855 ;
        RECT 108.505 155.625 108.795 155.855 ;
        RECT 108.965 155.810 109.255 155.855 ;
        RECT 109.410 155.810 109.730 155.870 ;
        RECT 108.965 155.670 109.730 155.810 ;
        RECT 108.965 155.625 109.255 155.670 ;
        RECT 105.360 155.470 105.500 155.610 ;
        RECT 108.580 155.470 108.720 155.625 ;
        RECT 105.360 155.330 108.720 155.470 ;
        RECT 109.040 155.130 109.180 155.625 ;
        RECT 109.410 155.610 109.730 155.670 ;
        RECT 113.090 155.810 113.410 155.870 ;
        RECT 116.325 155.810 116.615 155.855 ;
        RECT 113.090 155.670 116.615 155.810 ;
        RECT 113.090 155.610 113.410 155.670 ;
        RECT 116.325 155.625 116.615 155.670 ;
        RECT 117.690 155.270 118.010 155.530 ;
        RECT 108.580 154.990 109.180 155.130 ;
        RECT 106.650 154.790 106.970 154.850 ;
        RECT 108.580 154.790 108.720 154.990 ;
        RECT 104.900 154.650 108.720 154.790 ;
        RECT 110.345 154.790 110.635 154.835 ;
        RECT 110.790 154.790 111.110 154.850 ;
        RECT 110.345 154.650 111.110 154.790 ;
        RECT 103.445 154.605 103.735 154.650 ;
        RECT 103.890 154.590 104.210 154.650 ;
        RECT 106.650 154.590 106.970 154.650 ;
        RECT 110.345 154.605 110.635 154.650 ;
        RECT 110.790 154.590 111.110 154.650 ;
        RECT 14.580 153.970 127.740 154.450 ;
        RECT 23.865 153.770 24.155 153.815 ;
        RECT 27.530 153.770 27.850 153.830 ;
        RECT 23.865 153.630 27.850 153.770 ;
        RECT 23.865 153.585 24.155 153.630 ;
        RECT 27.530 153.570 27.850 153.630 ;
        RECT 70.310 153.770 70.630 153.830 ;
        RECT 72.165 153.770 72.455 153.815 ;
        RECT 70.310 153.630 72.455 153.770 ;
        RECT 70.310 153.570 70.630 153.630 ;
        RECT 72.165 153.585 72.455 153.630 ;
        RECT 73.530 153.570 73.850 153.830 ;
        RECT 98.830 153.770 99.150 153.830 ;
        RECT 84.890 153.630 99.150 153.770 ;
        RECT 33.940 153.430 34.230 153.475 ;
        RECT 36.720 153.430 37.010 153.475 ;
        RECT 38.580 153.430 38.870 153.475 ;
        RECT 54.210 153.430 54.530 153.490 ;
        RECT 33.940 153.290 38.870 153.430 ;
        RECT 33.940 153.245 34.230 153.290 ;
        RECT 36.720 153.245 37.010 153.290 ;
        RECT 38.580 153.245 38.870 153.290 ;
        RECT 42.340 153.290 54.530 153.430 ;
        RECT 21.090 152.890 21.410 153.150 ;
        RECT 21.565 153.090 21.855 153.135 ;
        RECT 22.010 153.090 22.330 153.150 ;
        RECT 21.565 152.950 22.330 153.090 ;
        RECT 21.565 152.905 21.855 152.950 ;
        RECT 22.010 152.890 22.330 152.950 ;
        RECT 37.190 152.890 37.510 153.150 ;
        RECT 37.650 153.090 37.970 153.150 ;
        RECT 37.650 152.950 42.020 153.090 ;
        RECT 37.650 152.890 37.970 152.950 ;
        RECT 33.940 152.750 34.230 152.795 ;
        RECT 36.730 152.750 37.050 152.810 ;
        RECT 41.880 152.795 42.020 152.950 ;
        RECT 39.045 152.750 39.335 152.795 ;
        RECT 33.940 152.610 36.475 152.750 ;
        RECT 33.940 152.565 34.230 152.610 ;
        RECT 32.080 152.410 32.370 152.455 ;
        RECT 33.510 152.410 33.830 152.470 ;
        RECT 36.260 152.455 36.475 152.610 ;
        RECT 36.730 152.610 39.335 152.750 ;
        RECT 36.730 152.550 37.050 152.610 ;
        RECT 39.045 152.565 39.335 152.610 ;
        RECT 40.885 152.565 41.175 152.795 ;
        RECT 41.345 152.565 41.635 152.795 ;
        RECT 41.805 152.565 42.095 152.795 ;
        RECT 35.340 152.410 35.630 152.455 ;
        RECT 32.080 152.270 35.630 152.410 ;
        RECT 32.080 152.225 32.370 152.270 ;
        RECT 33.510 152.210 33.830 152.270 ;
        RECT 35.340 152.225 35.630 152.270 ;
        RECT 36.260 152.410 36.550 152.455 ;
        RECT 38.120 152.410 38.410 152.455 ;
        RECT 36.260 152.270 38.410 152.410 ;
        RECT 36.260 152.225 36.550 152.270 ;
        RECT 38.120 152.225 38.410 152.270 ;
        RECT 22.025 152.070 22.315 152.115 ;
        RECT 22.470 152.070 22.790 152.130 ;
        RECT 22.025 151.930 22.790 152.070 ;
        RECT 22.025 151.885 22.315 151.930 ;
        RECT 22.470 151.870 22.790 151.930 ;
        RECT 30.075 152.070 30.365 152.115 ;
        RECT 31.210 152.070 31.530 152.130 ;
        RECT 30.075 151.930 31.530 152.070 ;
        RECT 30.075 151.885 30.365 151.930 ;
        RECT 31.210 151.870 31.530 151.930 ;
        RECT 34.890 152.070 35.210 152.130 ;
        RECT 39.505 152.070 39.795 152.115 ;
        RECT 34.890 151.930 39.795 152.070 ;
        RECT 40.960 152.070 41.100 152.565 ;
        RECT 41.420 152.410 41.560 152.565 ;
        RECT 42.340 152.410 42.480 153.290 ;
        RECT 54.210 153.230 54.530 153.290 ;
        RECT 62.460 153.430 62.750 153.475 ;
        RECT 65.240 153.430 65.530 153.475 ;
        RECT 67.100 153.430 67.390 153.475 ;
        RECT 62.460 153.290 67.390 153.430 ;
        RECT 62.460 153.245 62.750 153.290 ;
        RECT 65.240 153.245 65.530 153.290 ;
        RECT 67.100 153.245 67.390 153.290 ;
        RECT 69.850 153.430 70.170 153.490 ;
        RECT 84.890 153.430 85.030 153.630 ;
        RECT 98.830 153.570 99.150 153.630 ;
        RECT 102.970 153.770 103.290 153.830 ;
        RECT 103.445 153.770 103.735 153.815 ;
        RECT 109.870 153.770 110.190 153.830 ;
        RECT 102.970 153.630 103.735 153.770 ;
        RECT 102.970 153.570 103.290 153.630 ;
        RECT 103.445 153.585 103.735 153.630 ;
        RECT 107.200 153.630 110.190 153.770 ;
        RECT 69.850 153.290 85.030 153.430 ;
        RECT 90.520 153.430 90.810 153.475 ;
        RECT 93.300 153.430 93.590 153.475 ;
        RECT 95.160 153.430 95.450 153.475 ;
        RECT 90.520 153.290 95.450 153.430 ;
        RECT 98.920 153.430 99.060 153.570 ;
        RECT 105.270 153.430 105.590 153.490 ;
        RECT 98.920 153.290 105.590 153.430 ;
        RECT 69.850 153.230 70.170 153.290 ;
        RECT 90.520 153.245 90.810 153.290 ;
        RECT 93.300 153.245 93.590 153.290 ;
        RECT 95.160 153.245 95.450 153.290 ;
        RECT 105.270 153.230 105.590 153.290 ;
        RECT 64.330 153.090 64.650 153.150 ;
        RECT 69.390 153.090 69.710 153.150 ;
        RECT 73.990 153.090 74.310 153.150 ;
        RECT 74.465 153.090 74.755 153.135 ;
        RECT 64.330 152.950 69.160 153.090 ;
        RECT 64.330 152.890 64.650 152.950 ;
        RECT 42.725 152.750 43.015 152.795 ;
        RECT 44.550 152.750 44.870 152.810 ;
        RECT 42.725 152.610 44.870 152.750 ;
        RECT 42.725 152.565 43.015 152.610 ;
        RECT 44.550 152.550 44.870 152.610 ;
        RECT 50.990 152.750 51.310 152.810 ;
        RECT 56.970 152.750 57.290 152.810 ;
        RECT 50.990 152.610 57.290 152.750 ;
        RECT 50.990 152.550 51.310 152.610 ;
        RECT 56.970 152.550 57.290 152.610 ;
        RECT 62.460 152.750 62.750 152.795 ;
        RECT 62.460 152.610 64.995 152.750 ;
        RECT 62.460 152.565 62.750 152.610 ;
        RECT 43.170 152.410 43.490 152.470 ;
        RECT 64.780 152.455 64.995 152.610 ;
        RECT 65.710 152.550 66.030 152.810 ;
        RECT 67.565 152.750 67.855 152.795 ;
        RECT 68.470 152.750 68.790 152.810 ;
        RECT 67.565 152.610 68.790 152.750 ;
        RECT 69.020 152.750 69.160 152.950 ;
        RECT 69.390 152.950 73.760 153.090 ;
        RECT 69.390 152.890 69.710 152.950 ;
        RECT 70.770 152.750 71.090 152.810 ;
        RECT 69.020 152.610 71.090 152.750 ;
        RECT 67.565 152.565 67.855 152.610 ;
        RECT 68.470 152.550 68.790 152.610 ;
        RECT 70.770 152.550 71.090 152.610 ;
        RECT 71.245 152.565 71.535 152.795 ;
        RECT 71.690 152.750 72.010 152.810 ;
        RECT 73.085 152.750 73.375 152.795 ;
        RECT 71.690 152.610 73.375 152.750 ;
        RECT 73.620 152.750 73.760 152.950 ;
        RECT 73.990 152.950 74.755 153.090 ;
        RECT 73.990 152.890 74.310 152.950 ;
        RECT 74.465 152.905 74.755 152.950 ;
        RECT 91.930 153.090 92.250 153.150 ;
        RECT 91.930 152.950 93.540 153.090 ;
        RECT 91.930 152.890 92.250 152.950 ;
        RECT 74.925 152.750 75.215 152.795 ;
        RECT 73.620 152.610 75.215 152.750 ;
        RECT 41.420 152.270 43.490 152.410 ;
        RECT 43.170 152.210 43.490 152.270 ;
        RECT 57.445 152.410 57.735 152.455 ;
        RECT 60.600 152.410 60.890 152.455 ;
        RECT 63.860 152.410 64.150 152.455 ;
        RECT 57.445 152.270 64.150 152.410 ;
        RECT 57.445 152.225 57.735 152.270 ;
        RECT 60.600 152.225 60.890 152.270 ;
        RECT 63.860 152.225 64.150 152.270 ;
        RECT 64.780 152.410 65.070 152.455 ;
        RECT 66.640 152.410 66.930 152.455 ;
        RECT 64.780 152.270 66.930 152.410 ;
        RECT 71.320 152.410 71.460 152.565 ;
        RECT 71.690 152.550 72.010 152.610 ;
        RECT 73.085 152.565 73.375 152.610 ;
        RECT 74.925 152.565 75.215 152.610 ;
        RECT 90.520 152.750 90.810 152.795 ;
        RECT 93.400 152.750 93.540 152.950 ;
        RECT 93.770 152.890 94.090 153.150 ;
        RECT 104.350 152.890 104.670 153.150 ;
        RECT 105.360 153.090 105.500 153.230 ;
        RECT 107.200 153.090 107.340 153.630 ;
        RECT 109.870 153.570 110.190 153.630 ;
        RECT 108.030 153.430 108.350 153.490 ;
        RECT 114.470 153.430 114.790 153.490 ;
        RECT 108.030 153.290 114.790 153.430 ;
        RECT 108.030 153.230 108.350 153.290 ;
        RECT 114.470 153.230 114.790 153.290 ;
        RECT 105.360 152.950 107.340 153.090 ;
        RECT 95.625 152.750 95.915 152.795 ;
        RECT 90.520 152.610 93.055 152.750 ;
        RECT 93.400 152.610 95.915 152.750 ;
        RECT 90.520 152.565 90.810 152.610 ;
        RECT 72.150 152.410 72.470 152.470 ;
        RECT 73.530 152.410 73.850 152.470 ;
        RECT 87.790 152.410 88.110 152.470 ;
        RECT 92.840 152.455 93.055 152.610 ;
        RECT 95.625 152.565 95.915 152.610 ;
        RECT 103.445 152.750 103.735 152.795 ;
        RECT 103.445 152.610 106.420 152.750 ;
        RECT 103.445 152.565 103.735 152.610 ;
        RECT 71.320 152.270 73.850 152.410 ;
        RECT 64.780 152.225 65.070 152.270 ;
        RECT 66.640 152.225 66.930 152.270 ;
        RECT 72.150 152.210 72.470 152.270 ;
        RECT 73.530 152.210 73.850 152.270 ;
        RECT 74.540 152.270 88.110 152.410 ;
        RECT 41.790 152.070 42.110 152.130 ;
        RECT 50.530 152.070 50.850 152.130 ;
        RECT 58.810 152.115 59.130 152.130 ;
        RECT 40.960 151.930 50.850 152.070 ;
        RECT 34.890 151.870 35.210 151.930 ;
        RECT 39.505 151.885 39.795 151.930 ;
        RECT 41.790 151.870 42.110 151.930 ;
        RECT 50.530 151.870 50.850 151.930 ;
        RECT 58.595 151.885 59.130 152.115 ;
        RECT 58.810 151.870 59.130 151.885 ;
        RECT 70.310 152.070 70.630 152.130 ;
        RECT 74.540 152.070 74.680 152.270 ;
        RECT 87.790 152.210 88.110 152.270 ;
        RECT 88.660 152.410 88.950 152.455 ;
        RECT 91.920 152.410 92.210 152.455 ;
        RECT 92.840 152.410 93.130 152.455 ;
        RECT 94.700 152.410 94.990 152.455 ;
        RECT 88.660 152.270 92.620 152.410 ;
        RECT 88.660 152.225 88.950 152.270 ;
        RECT 91.920 152.225 92.210 152.270 ;
        RECT 70.310 151.930 74.680 152.070 ;
        RECT 70.310 151.870 70.630 151.930 ;
        RECT 74.910 151.870 75.230 152.130 ;
        RECT 86.410 152.115 86.730 152.130 ;
        RECT 86.410 151.885 86.945 152.115 ;
        RECT 92.480 152.070 92.620 152.270 ;
        RECT 92.840 152.270 94.990 152.410 ;
        RECT 92.840 152.225 93.130 152.270 ;
        RECT 94.700 152.225 94.990 152.270 ;
        RECT 104.810 152.210 105.130 152.470 ;
        RECT 106.280 152.410 106.420 152.610 ;
        RECT 106.650 152.550 106.970 152.810 ;
        RECT 107.200 152.795 107.340 152.950 ;
        RECT 109.870 153.090 110.190 153.150 ;
        RECT 116.310 153.090 116.630 153.150 ;
        RECT 109.870 152.950 111.020 153.090 ;
        RECT 109.870 152.890 110.190 152.950 ;
        RECT 107.125 152.565 107.415 152.795 ;
        RECT 107.570 152.550 107.890 152.810 ;
        RECT 108.490 152.550 108.810 152.810 ;
        RECT 109.410 152.750 109.730 152.810 ;
        RECT 110.880 152.795 111.020 152.950 ;
        RECT 111.340 152.950 116.630 153.090 ;
        RECT 111.340 152.795 111.480 152.950 ;
        RECT 116.310 152.890 116.630 152.950 ;
        RECT 110.345 152.750 110.635 152.795 ;
        RECT 109.410 152.610 110.635 152.750 ;
        RECT 109.410 152.550 109.730 152.610 ;
        RECT 110.345 152.565 110.635 152.610 ;
        RECT 110.805 152.565 111.095 152.795 ;
        RECT 111.265 152.565 111.555 152.795 ;
        RECT 112.185 152.750 112.475 152.795 ;
        RECT 119.530 152.750 119.850 152.810 ;
        RECT 111.800 152.610 112.475 152.750 ;
        RECT 108.965 152.410 109.255 152.455 ;
        RECT 106.280 152.270 109.255 152.410 ;
        RECT 108.965 152.225 109.255 152.270 ;
        RECT 93.770 152.070 94.090 152.130 ;
        RECT 92.480 151.930 94.090 152.070 ;
        RECT 86.410 151.870 86.730 151.885 ;
        RECT 93.770 151.870 94.090 151.930 ;
        RECT 101.590 152.070 101.910 152.130 ;
        RECT 102.525 152.070 102.815 152.115 ;
        RECT 101.590 151.930 102.815 152.070 ;
        RECT 101.590 151.870 101.910 151.930 ;
        RECT 102.525 151.885 102.815 151.930 ;
        RECT 105.270 151.870 105.590 152.130 ;
        RECT 108.490 152.070 108.810 152.130 ;
        RECT 111.800 152.070 111.940 152.610 ;
        RECT 112.185 152.565 112.475 152.610 ;
        RECT 112.720 152.610 119.850 152.750 ;
        RECT 108.490 151.930 111.940 152.070 ;
        RECT 112.170 152.070 112.490 152.130 ;
        RECT 112.720 152.070 112.860 152.610 ;
        RECT 119.530 152.550 119.850 152.610 ;
        RECT 120.465 152.565 120.755 152.795 ;
        RECT 115.850 152.410 116.170 152.470 ;
        RECT 120.540 152.410 120.680 152.565 ;
        RECT 115.850 152.270 120.680 152.410 ;
        RECT 115.850 152.210 116.170 152.270 ;
        RECT 112.170 151.930 112.860 152.070 ;
        RECT 118.150 152.070 118.470 152.130 ;
        RECT 119.085 152.070 119.375 152.115 ;
        RECT 118.150 151.930 119.375 152.070 ;
        RECT 108.490 151.870 108.810 151.930 ;
        RECT 112.170 151.870 112.490 151.930 ;
        RECT 118.150 151.870 118.470 151.930 ;
        RECT 119.085 151.885 119.375 151.930 ;
        RECT 121.385 152.070 121.675 152.115 ;
        RECT 123.210 152.070 123.530 152.130 ;
        RECT 121.385 151.930 123.530 152.070 ;
        RECT 121.385 151.885 121.675 151.930 ;
        RECT 123.210 151.870 123.530 151.930 ;
        RECT 14.580 151.250 127.740 151.730 ;
        RECT 33.510 150.850 33.830 151.110 ;
        RECT 36.745 151.050 37.035 151.095 ;
        RECT 37.190 151.050 37.510 151.110 ;
        RECT 36.745 150.910 37.510 151.050 ;
        RECT 36.745 150.865 37.035 150.910 ;
        RECT 37.190 150.850 37.510 150.910 ;
        RECT 60.665 150.865 60.955 151.095 ;
        RECT 61.110 151.050 61.430 151.110 ;
        RECT 61.585 151.050 61.875 151.095 ;
        RECT 61.110 150.910 61.875 151.050 ;
        RECT 18.740 150.710 19.030 150.755 ;
        RECT 20.170 150.710 20.490 150.770 ;
        RECT 22.000 150.710 22.290 150.755 ;
        RECT 18.740 150.570 22.290 150.710 ;
        RECT 18.740 150.525 19.030 150.570 ;
        RECT 20.170 150.510 20.490 150.570 ;
        RECT 22.000 150.525 22.290 150.570 ;
        RECT 22.920 150.710 23.210 150.755 ;
        RECT 24.780 150.710 25.070 150.755 ;
        RECT 22.920 150.570 25.070 150.710 ;
        RECT 22.920 150.525 23.210 150.570 ;
        RECT 24.780 150.525 25.070 150.570 ;
        RECT 31.210 150.710 31.530 150.770 ;
        RECT 58.365 150.710 58.655 150.755 ;
        RECT 31.210 150.570 43.860 150.710 ;
        RECT 20.600 150.370 20.890 150.415 ;
        RECT 22.920 150.370 23.135 150.525 ;
        RECT 31.210 150.510 31.530 150.570 ;
        RECT 20.600 150.230 23.135 150.370 ;
        RECT 29.830 150.370 30.150 150.430 ;
        RECT 33.065 150.370 33.355 150.415 ;
        RECT 29.830 150.230 33.355 150.370 ;
        RECT 20.600 150.185 20.890 150.230 ;
        RECT 29.830 150.170 30.150 150.230 ;
        RECT 33.065 150.185 33.355 150.230 ;
        RECT 35.810 150.170 36.130 150.430 ;
        RECT 41.790 150.370 42.110 150.430 ;
        RECT 42.725 150.370 43.015 150.415 ;
        RECT 41.790 150.230 43.015 150.370 ;
        RECT 41.790 150.170 42.110 150.230 ;
        RECT 42.725 150.185 43.015 150.230 ;
        RECT 43.170 150.170 43.490 150.430 ;
        RECT 43.720 150.415 43.860 150.570 ;
        RECT 53.840 150.570 58.655 150.710 ;
        RECT 53.840 150.430 53.980 150.570 ;
        RECT 58.365 150.525 58.655 150.570 ;
        RECT 43.645 150.185 43.935 150.415 ;
        RECT 44.565 150.370 44.855 150.415 ;
        RECT 45.010 150.370 45.330 150.430 ;
        RECT 44.565 150.230 45.330 150.370 ;
        RECT 44.565 150.185 44.855 150.230 ;
        RECT 45.010 150.170 45.330 150.230 ;
        RECT 48.705 150.185 48.995 150.415 ;
        RECT 16.735 150.030 17.025 150.075 ;
        RECT 22.470 150.030 22.790 150.090 ;
        RECT 16.735 149.890 22.790 150.030 ;
        RECT 16.735 149.845 17.025 149.890 ;
        RECT 22.470 149.830 22.790 149.890 ;
        RECT 23.865 150.030 24.155 150.075 ;
        RECT 24.770 150.030 25.090 150.090 ;
        RECT 23.865 149.890 25.090 150.030 ;
        RECT 23.865 149.845 24.155 149.890 ;
        RECT 24.770 149.830 25.090 149.890 ;
        RECT 25.705 150.030 25.995 150.075 ;
        RECT 36.270 150.030 36.590 150.090 ;
        RECT 25.705 149.890 36.590 150.030 ;
        RECT 48.780 150.030 48.920 150.185 ;
        RECT 49.610 150.170 49.930 150.430 ;
        RECT 50.070 150.170 50.390 150.430 ;
        RECT 52.845 150.185 53.135 150.415 ;
        RECT 50.530 150.030 50.850 150.090 ;
        RECT 48.780 149.890 50.850 150.030 ;
        RECT 52.920 150.030 53.060 150.185 ;
        RECT 53.290 150.170 53.610 150.430 ;
        RECT 53.750 150.170 54.070 150.430 ;
        RECT 54.685 150.370 54.975 150.415 ;
        RECT 56.510 150.370 56.830 150.430 ;
        RECT 54.685 150.230 56.830 150.370 ;
        RECT 54.685 150.185 54.975 150.230 ;
        RECT 56.510 150.170 56.830 150.230 ;
        RECT 58.810 150.170 59.130 150.430 ;
        RECT 60.740 150.370 60.880 150.865 ;
        RECT 61.110 150.850 61.430 150.910 ;
        RECT 61.585 150.865 61.875 150.910 ;
        RECT 64.805 151.050 65.095 151.095 ;
        RECT 65.710 151.050 66.030 151.110 ;
        RECT 64.805 150.910 66.030 151.050 ;
        RECT 64.805 150.865 65.095 150.910 ;
        RECT 65.710 150.850 66.030 150.910 ;
        RECT 68.485 151.050 68.775 151.095 ;
        RECT 85.965 151.050 86.255 151.095 ;
        RECT 86.410 151.050 86.730 151.110 ;
        RECT 88.265 151.050 88.555 151.095 ;
        RECT 92.865 151.050 93.155 151.095 ;
        RECT 93.310 151.050 93.630 151.110 ;
        RECT 68.485 150.910 71.460 151.050 ;
        RECT 68.485 150.865 68.775 150.910 ;
        RECT 62.505 150.370 62.795 150.415 ;
        RECT 60.740 150.230 62.795 150.370 ;
        RECT 62.505 150.185 62.795 150.230 ;
        RECT 63.870 150.170 64.190 150.430 ;
        RECT 67.565 150.370 67.855 150.415 ;
        RECT 69.390 150.370 69.710 150.430 ;
        RECT 67.565 150.230 69.710 150.370 ;
        RECT 67.565 150.185 67.855 150.230 ;
        RECT 69.390 150.170 69.710 150.230 ;
        RECT 70.770 150.170 71.090 150.430 ;
        RECT 54.210 150.030 54.530 150.090 ;
        RECT 52.920 149.890 54.530 150.030 ;
        RECT 25.705 149.845 25.995 149.890 ;
        RECT 36.270 149.830 36.590 149.890 ;
        RECT 50.530 149.830 50.850 149.890 ;
        RECT 54.210 149.830 54.530 149.890 ;
        RECT 57.905 150.030 58.195 150.075 ;
        RECT 65.710 150.030 66.030 150.090 ;
        RECT 57.905 149.890 65.020 150.030 ;
        RECT 57.905 149.845 58.195 149.890 ;
        RECT 64.880 149.750 65.020 149.890 ;
        RECT 65.710 149.890 71.000 150.030 ;
        RECT 65.710 149.830 66.030 149.890 ;
        RECT 20.600 149.690 20.890 149.735 ;
        RECT 23.380 149.690 23.670 149.735 ;
        RECT 25.240 149.690 25.530 149.735 ;
        RECT 20.600 149.550 25.530 149.690 ;
        RECT 20.600 149.505 20.890 149.550 ;
        RECT 23.380 149.505 23.670 149.550 ;
        RECT 25.240 149.505 25.530 149.550 ;
        RECT 51.005 149.690 51.295 149.735 ;
        RECT 60.190 149.690 60.510 149.750 ;
        RECT 51.005 149.550 60.510 149.690 ;
        RECT 51.005 149.505 51.295 149.550 ;
        RECT 60.190 149.490 60.510 149.550 ;
        RECT 64.790 149.690 65.110 149.750 ;
        RECT 70.860 149.690 71.000 149.890 ;
        RECT 71.320 149.690 71.460 150.910 ;
        RECT 85.965 150.910 87.100 151.050 ;
        RECT 85.965 150.865 86.255 150.910 ;
        RECT 86.410 150.850 86.730 150.910 ;
        RECT 73.085 150.710 73.375 150.755 ;
        RECT 74.910 150.710 75.230 150.770 ;
        RECT 75.385 150.710 75.675 150.755 ;
        RECT 73.085 150.570 75.675 150.710 ;
        RECT 73.085 150.525 73.375 150.570 ;
        RECT 74.910 150.510 75.230 150.570 ;
        RECT 75.385 150.525 75.675 150.570 ;
        RECT 77.225 150.710 77.515 150.755 ;
        RECT 77.225 150.570 85.260 150.710 ;
        RECT 77.225 150.525 77.515 150.570 ;
        RECT 75.830 150.370 76.150 150.430 ;
        RECT 78.605 150.370 78.895 150.415 ;
        RECT 75.830 150.230 78.895 150.370 ;
        RECT 75.830 150.170 76.150 150.230 ;
        RECT 78.605 150.185 78.895 150.230 ;
        RECT 79.970 150.170 80.290 150.430 ;
        RECT 85.120 150.090 85.260 150.570 ;
        RECT 85.950 150.370 86.270 150.430 ;
        RECT 86.425 150.370 86.715 150.415 ;
        RECT 85.950 150.230 86.715 150.370 ;
        RECT 85.950 150.170 86.270 150.230 ;
        RECT 86.425 150.185 86.715 150.230 ;
        RECT 79.510 149.830 79.830 150.090 ;
        RECT 85.030 149.830 85.350 150.090 ;
        RECT 78.130 149.690 78.450 149.750 ;
        RECT 64.790 149.550 70.540 149.690 ;
        RECT 70.860 149.550 78.450 149.690 ;
        RECT 86.960 149.690 87.100 150.910 ;
        RECT 88.265 150.910 92.160 151.050 ;
        RECT 88.265 150.865 88.555 150.910 ;
        RECT 92.020 150.535 92.160 150.910 ;
        RECT 92.865 150.910 93.630 151.050 ;
        RECT 92.865 150.865 93.155 150.910 ;
        RECT 93.310 150.850 93.630 150.910 ;
        RECT 93.770 150.850 94.090 151.110 ;
        RECT 104.810 151.050 105.130 151.110 ;
        RECT 107.125 151.050 107.415 151.095 ;
        RECT 94.320 150.910 104.580 151.050 ;
        RECT 90.565 150.185 90.855 150.415 ;
        RECT 91.945 150.305 92.235 150.535 ;
        RECT 94.320 150.415 94.460 150.910 ;
        RECT 95.610 150.710 95.930 150.770 ;
        RECT 98.025 150.710 98.315 150.755 ;
        RECT 101.265 150.710 101.915 150.755 ;
        RECT 95.610 150.570 101.915 150.710 ;
        RECT 95.610 150.510 95.930 150.570 ;
        RECT 98.025 150.525 98.615 150.570 ;
        RECT 101.265 150.525 101.915 150.570 ;
        RECT 103.430 150.710 103.750 150.770 ;
        RECT 103.905 150.710 104.195 150.755 ;
        RECT 103.430 150.570 104.195 150.710 ;
        RECT 104.440 150.710 104.580 150.910 ;
        RECT 104.810 150.910 107.415 151.050 ;
        RECT 104.810 150.850 105.130 150.910 ;
        RECT 107.125 150.865 107.415 150.910 ;
        RECT 116.770 150.710 117.090 150.770 ;
        RECT 104.440 150.570 117.090 150.710 ;
        RECT 94.245 150.370 94.535 150.415 ;
        RECT 92.480 150.230 94.535 150.370 ;
        RECT 90.640 150.030 90.780 150.185 ;
        RECT 92.480 150.030 92.620 150.230 ;
        RECT 94.245 150.185 94.535 150.230 ;
        RECT 98.325 150.210 98.615 150.525 ;
        RECT 103.430 150.510 103.750 150.570 ;
        RECT 103.905 150.525 104.195 150.570 ;
        RECT 116.770 150.510 117.090 150.570 ;
        RECT 117.345 150.710 117.635 150.755 ;
        RECT 118.150 150.710 118.470 150.770 ;
        RECT 120.585 150.710 121.235 150.755 ;
        RECT 117.345 150.570 121.235 150.710 ;
        RECT 117.345 150.525 117.935 150.570 ;
        RECT 99.405 150.370 99.695 150.415 ;
        RECT 102.985 150.370 103.275 150.415 ;
        RECT 104.820 150.370 105.110 150.415 ;
        RECT 99.405 150.230 105.110 150.370 ;
        RECT 99.405 150.185 99.695 150.230 ;
        RECT 102.985 150.185 103.275 150.230 ;
        RECT 104.820 150.185 105.110 150.230 ;
        RECT 108.030 150.370 108.350 150.430 ;
        RECT 108.505 150.370 108.795 150.415 ;
        RECT 108.030 150.230 108.795 150.370 ;
        RECT 108.030 150.170 108.350 150.230 ;
        RECT 108.505 150.185 108.795 150.230 ;
        RECT 108.965 150.185 109.255 150.415 ;
        RECT 109.425 150.185 109.715 150.415 ;
        RECT 109.870 150.370 110.190 150.430 ;
        RECT 110.345 150.370 110.635 150.415 ;
        RECT 109.870 150.230 110.635 150.370 ;
        RECT 105.285 150.030 105.575 150.075 ;
        RECT 90.640 149.890 92.620 150.030 ;
        RECT 94.320 149.890 105.575 150.030 ;
        RECT 94.320 149.750 94.460 149.890 ;
        RECT 105.285 149.845 105.575 149.890 ;
        RECT 107.570 150.030 107.890 150.090 ;
        RECT 109.040 150.030 109.180 150.185 ;
        RECT 107.570 149.890 109.180 150.030 ;
        RECT 109.500 150.030 109.640 150.185 ;
        RECT 109.870 150.170 110.190 150.230 ;
        RECT 110.345 150.185 110.635 150.230 ;
        RECT 117.645 150.210 117.935 150.525 ;
        RECT 118.150 150.510 118.470 150.570 ;
        RECT 120.585 150.525 121.235 150.570 ;
        RECT 123.210 150.510 123.530 150.770 ;
        RECT 118.725 150.370 119.015 150.415 ;
        RECT 122.305 150.370 122.595 150.415 ;
        RECT 124.140 150.370 124.430 150.415 ;
        RECT 118.725 150.230 124.430 150.370 ;
        RECT 118.725 150.185 119.015 150.230 ;
        RECT 122.305 150.185 122.595 150.230 ;
        RECT 124.140 150.185 124.430 150.230 ;
        RECT 111.265 150.030 111.555 150.075 ;
        RECT 115.865 150.030 116.155 150.075 ;
        RECT 109.500 149.890 116.155 150.030 ;
        RECT 107.570 149.830 107.890 149.890 ;
        RECT 93.770 149.690 94.090 149.750 ;
        RECT 86.960 149.550 94.090 149.690 ;
        RECT 64.790 149.490 65.110 149.550 ;
        RECT 40.870 149.350 41.190 149.410 ;
        RECT 41.345 149.350 41.635 149.395 ;
        RECT 40.870 149.210 41.635 149.350 ;
        RECT 40.870 149.150 41.190 149.210 ;
        RECT 41.345 149.165 41.635 149.210 ;
        RECT 44.090 149.350 44.410 149.410 ;
        RECT 48.705 149.350 48.995 149.395 ;
        RECT 44.090 149.210 48.995 149.350 ;
        RECT 44.090 149.150 44.410 149.210 ;
        RECT 48.705 149.165 48.995 149.210 ;
        RECT 51.450 149.150 51.770 149.410 ;
        RECT 65.250 149.350 65.570 149.410 ;
        RECT 69.865 149.350 70.155 149.395 ;
        RECT 65.250 149.210 70.155 149.350 ;
        RECT 70.400 149.350 70.540 149.550 ;
        RECT 78.130 149.490 78.450 149.550 ;
        RECT 93.770 149.490 94.090 149.550 ;
        RECT 94.230 149.490 94.550 149.750 ;
        RECT 99.405 149.690 99.695 149.735 ;
        RECT 102.525 149.690 102.815 149.735 ;
        RECT 104.415 149.690 104.705 149.735 ;
        RECT 99.405 149.550 104.705 149.690 ;
        RECT 109.040 149.690 109.180 149.890 ;
        RECT 111.265 149.845 111.555 149.890 ;
        RECT 115.865 149.845 116.155 149.890 ;
        RECT 124.605 150.030 124.895 150.075 ;
        RECT 125.970 150.030 126.290 150.090 ;
        RECT 124.605 149.890 126.290 150.030 ;
        RECT 124.605 149.845 124.895 149.890 ;
        RECT 125.970 149.830 126.290 149.890 ;
        RECT 111.710 149.690 112.030 149.750 ;
        RECT 109.040 149.550 112.030 149.690 ;
        RECT 99.405 149.505 99.695 149.550 ;
        RECT 102.525 149.505 102.815 149.550 ;
        RECT 104.415 149.505 104.705 149.550 ;
        RECT 111.710 149.490 112.030 149.550 ;
        RECT 118.725 149.690 119.015 149.735 ;
        RECT 121.845 149.690 122.135 149.735 ;
        RECT 123.735 149.690 124.025 149.735 ;
        RECT 118.725 149.550 124.025 149.690 ;
        RECT 118.725 149.505 119.015 149.550 ;
        RECT 121.845 149.505 122.135 149.550 ;
        RECT 123.735 149.505 124.025 149.550 ;
        RECT 71.705 149.350 71.995 149.395 ;
        RECT 70.400 149.210 71.995 149.350 ;
        RECT 65.250 149.150 65.570 149.210 ;
        RECT 69.865 149.165 70.155 149.210 ;
        RECT 71.705 149.165 71.995 149.210 ;
        RECT 75.830 149.350 76.150 149.410 ;
        RECT 77.685 149.350 77.975 149.395 ;
        RECT 75.830 149.210 77.975 149.350 ;
        RECT 75.830 149.150 76.150 149.210 ;
        RECT 77.685 149.165 77.975 149.210 ;
        RECT 79.985 149.350 80.275 149.395 ;
        RECT 81.810 149.350 82.130 149.410 ;
        RECT 79.985 149.210 82.130 149.350 ;
        RECT 79.985 149.165 80.275 149.210 ;
        RECT 81.810 149.150 82.130 149.210 ;
        RECT 90.105 149.350 90.395 149.395 ;
        RECT 90.550 149.350 90.870 149.410 ;
        RECT 90.105 149.210 90.870 149.350 ;
        RECT 90.105 149.165 90.395 149.210 ;
        RECT 90.550 149.150 90.870 149.210 ;
        RECT 96.530 149.150 96.850 149.410 ;
        RECT 114.010 149.150 114.330 149.410 ;
        RECT 14.580 148.530 127.740 149.010 ;
        RECT 24.770 148.130 25.090 148.390 ;
        RECT 35.810 148.330 36.130 148.390 ;
        RECT 48.705 148.330 48.995 148.375 ;
        RECT 49.150 148.330 49.470 148.390 ;
        RECT 35.810 148.190 42.940 148.330 ;
        RECT 35.810 148.130 36.130 148.190 ;
        RECT 23.865 147.805 24.155 148.035 ;
        RECT 28.450 147.990 28.770 148.050 ;
        RECT 28.450 147.850 34.660 147.990 ;
        RECT 21.090 147.450 21.410 147.710 ;
        RECT 23.940 147.310 24.080 147.805 ;
        RECT 28.450 147.790 28.770 147.850 ;
        RECT 32.605 147.650 32.895 147.695 ;
        RECT 33.970 147.650 34.290 147.710 ;
        RECT 26.240 147.510 31.900 147.650 ;
        RECT 25.705 147.310 25.995 147.355 ;
        RECT 23.940 147.170 25.995 147.310 ;
        RECT 25.705 147.125 25.995 147.170 ;
        RECT 22.025 146.970 22.315 147.015 ;
        RECT 22.930 146.970 23.250 147.030 ;
        RECT 26.240 146.970 26.380 147.510 ;
        RECT 28.005 147.310 28.295 147.355 ;
        RECT 28.005 147.170 30.060 147.310 ;
        RECT 28.005 147.125 28.295 147.170 ;
        RECT 22.025 146.830 26.380 146.970 ;
        RECT 22.025 146.785 22.315 146.830 ;
        RECT 22.930 146.770 23.250 146.830 ;
        RECT 21.565 146.630 21.855 146.675 ;
        RECT 22.470 146.630 22.790 146.690 ;
        RECT 28.450 146.630 28.770 146.690 ;
        RECT 21.565 146.490 28.770 146.630 ;
        RECT 21.565 146.445 21.855 146.490 ;
        RECT 22.470 146.430 22.790 146.490 ;
        RECT 28.450 146.430 28.770 146.490 ;
        RECT 28.910 146.430 29.230 146.690 ;
        RECT 29.385 146.630 29.675 146.675 ;
        RECT 29.920 146.630 30.060 147.170 ;
        RECT 31.210 147.110 31.530 147.370 ;
        RECT 31.760 147.015 31.900 147.510 ;
        RECT 32.605 147.510 34.290 147.650 ;
        RECT 34.520 147.650 34.660 147.850 ;
        RECT 36.820 147.850 42.020 147.990 ;
        RECT 36.820 147.650 36.960 147.850 ;
        RECT 34.520 147.510 36.960 147.650 ;
        RECT 37.280 147.510 41.560 147.650 ;
        RECT 32.605 147.465 32.895 147.510 ;
        RECT 33.970 147.450 34.290 147.510 ;
        RECT 35.810 147.110 36.130 147.370 ;
        RECT 37.280 147.355 37.420 147.510 ;
        RECT 41.420 147.355 41.560 147.510 ;
        RECT 41.880 147.355 42.020 147.850 ;
        RECT 42.800 147.355 42.940 148.190 ;
        RECT 48.705 148.190 49.470 148.330 ;
        RECT 48.705 148.145 48.995 148.190 ;
        RECT 49.150 148.130 49.470 148.190 ;
        RECT 50.530 148.330 50.850 148.390 ;
        RECT 53.305 148.330 53.595 148.375 ;
        RECT 50.530 148.190 53.595 148.330 ;
        RECT 50.530 148.130 50.850 148.190 ;
        RECT 53.305 148.145 53.595 148.190 ;
        RECT 54.670 148.330 54.990 148.390 ;
        RECT 73.530 148.330 73.850 148.390 ;
        RECT 54.670 148.190 73.850 148.330 ;
        RECT 54.670 148.130 54.990 148.190 ;
        RECT 73.530 148.130 73.850 148.190 ;
        RECT 79.970 148.130 80.290 148.390 ;
        RECT 85.030 148.330 85.350 148.390 ;
        RECT 85.030 148.190 95.380 148.330 ;
        RECT 85.030 148.130 85.350 148.190 ;
        RECT 49.625 147.990 49.915 148.035 ;
        RECT 56.970 147.990 57.290 148.050 ;
        RECT 78.130 147.990 78.450 148.050 ;
        RECT 83.190 147.990 83.510 148.050 ;
        RECT 49.625 147.850 57.290 147.990 ;
        RECT 49.625 147.805 49.915 147.850 ;
        RECT 56.970 147.790 57.290 147.850 ;
        RECT 57.520 147.850 66.400 147.990 ;
        RECT 48.245 147.650 48.535 147.695 ;
        RECT 52.370 147.650 52.690 147.710 ;
        RECT 48.245 147.510 52.690 147.650 ;
        RECT 48.245 147.465 48.535 147.510 ;
        RECT 52.370 147.450 52.690 147.510 ;
        RECT 53.290 147.650 53.610 147.710 ;
        RECT 57.520 147.650 57.660 147.850 ;
        RECT 53.290 147.510 57.660 147.650 ;
        RECT 60.665 147.650 60.955 147.695 ;
        RECT 64.790 147.650 65.110 147.710 ;
        RECT 60.665 147.510 65.110 147.650 ;
        RECT 53.290 147.450 53.610 147.510 ;
        RECT 36.745 147.125 37.035 147.355 ;
        RECT 37.205 147.125 37.495 147.355 ;
        RECT 37.665 147.310 37.955 147.355 ;
        RECT 40.885 147.310 41.175 147.355 ;
        RECT 37.665 147.170 41.175 147.310 ;
        RECT 37.665 147.125 37.955 147.170 ;
        RECT 40.885 147.125 41.175 147.170 ;
        RECT 41.345 147.125 41.635 147.355 ;
        RECT 41.805 147.125 42.095 147.355 ;
        RECT 42.725 147.310 43.015 147.355 ;
        RECT 44.550 147.310 44.870 147.370 ;
        RECT 42.725 147.170 44.870 147.310 ;
        RECT 42.725 147.125 43.015 147.170 ;
        RECT 31.685 146.970 31.975 147.015 ;
        RECT 36.820 146.970 36.960 147.125 ;
        RECT 39.505 146.970 39.795 147.015 ;
        RECT 31.685 146.830 36.960 146.970 ;
        RECT 37.740 146.830 39.795 146.970 ;
        RECT 31.685 146.785 31.975 146.830 ;
        RECT 29.385 146.490 30.060 146.630 ;
        RECT 36.730 146.630 37.050 146.690 ;
        RECT 37.740 146.630 37.880 146.830 ;
        RECT 39.505 146.785 39.795 146.830 ;
        RECT 36.730 146.490 37.880 146.630 ;
        RECT 38.570 146.630 38.890 146.690 ;
        RECT 39.045 146.630 39.335 146.675 ;
        RECT 38.570 146.490 39.335 146.630 ;
        RECT 40.960 146.630 41.100 147.125 ;
        RECT 41.420 146.970 41.560 147.125 ;
        RECT 44.550 147.110 44.870 147.170 ;
        RECT 48.690 147.110 49.010 147.370 ;
        RECT 51.910 147.110 52.230 147.370 ;
        RECT 54.670 147.110 54.990 147.370 ;
        RECT 55.220 147.355 55.360 147.510 ;
        RECT 60.665 147.465 60.955 147.510 ;
        RECT 64.790 147.450 65.110 147.510 ;
        RECT 55.145 147.125 55.435 147.355 ;
        RECT 55.605 147.125 55.895 147.355 ;
        RECT 56.510 147.310 56.830 147.370 ;
        RECT 65.710 147.310 66.030 147.370 ;
        RECT 56.510 147.170 66.030 147.310 ;
        RECT 66.260 147.310 66.400 147.850 ;
        RECT 76.380 147.850 83.510 147.990 ;
        RECT 70.770 147.650 71.090 147.710 ;
        RECT 70.770 147.510 72.840 147.650 ;
        RECT 70.770 147.450 71.090 147.510 ;
        RECT 66.260 147.170 71.230 147.310 ;
        RECT 43.170 146.970 43.490 147.030 ;
        RECT 41.420 146.830 43.490 146.970 ;
        RECT 43.170 146.770 43.490 146.830 ;
        RECT 47.325 146.970 47.615 147.015 ;
        RECT 51.450 146.970 51.770 147.030 ;
        RECT 47.325 146.830 51.770 146.970 ;
        RECT 55.680 146.970 55.820 147.125 ;
        RECT 56.510 147.110 56.830 147.170 ;
        RECT 65.710 147.110 66.030 147.170 ;
        RECT 58.810 146.970 59.130 147.030 ;
        RECT 61.125 146.970 61.415 147.015 ;
        RECT 55.680 146.830 61.415 146.970 ;
        RECT 71.090 146.970 71.230 147.170 ;
        RECT 72.150 147.110 72.470 147.370 ;
        RECT 72.700 147.355 72.840 147.510 ;
        RECT 76.380 147.355 76.520 147.850 ;
        RECT 78.130 147.790 78.450 147.850 ;
        RECT 83.190 147.790 83.510 147.850 ;
        RECT 89.140 147.990 89.430 148.035 ;
        RECT 91.920 147.990 92.210 148.035 ;
        RECT 93.780 147.990 94.070 148.035 ;
        RECT 89.140 147.850 94.070 147.990 ;
        RECT 95.240 147.990 95.380 148.190 ;
        RECT 95.610 148.130 95.930 148.390 ;
        RECT 96.530 148.330 96.850 148.390 ;
        RECT 102.985 148.330 103.275 148.375 ;
        RECT 103.430 148.330 103.750 148.390 ;
        RECT 96.530 148.190 100.900 148.330 ;
        RECT 96.530 148.130 96.850 148.190 ;
        RECT 95.240 147.850 97.220 147.990 ;
        RECT 89.140 147.805 89.430 147.850 ;
        RECT 91.920 147.805 92.210 147.850 ;
        RECT 93.780 147.805 94.070 147.850 ;
        RECT 86.410 147.650 86.730 147.710 ;
        RECT 77.300 147.510 86.730 147.650 ;
        RECT 77.300 147.355 77.440 147.510 ;
        RECT 86.410 147.450 86.730 147.510 ;
        RECT 91.010 147.650 91.330 147.710 ;
        RECT 97.080 147.695 97.220 147.850 ;
        RECT 100.225 147.805 100.515 148.035 ;
        RECT 100.760 147.990 100.900 148.190 ;
        RECT 102.985 148.190 103.750 148.330 ;
        RECT 102.985 148.145 103.275 148.190 ;
        RECT 103.430 148.130 103.750 148.190 ;
        RECT 103.905 148.330 104.195 148.375 ;
        RECT 104.350 148.330 104.670 148.390 ;
        RECT 103.905 148.190 104.670 148.330 ;
        RECT 103.905 148.145 104.195 148.190 ;
        RECT 104.350 148.130 104.670 148.190 ;
        RECT 106.190 148.130 106.510 148.390 ;
        RECT 115.850 148.130 116.170 148.390 ;
        RECT 120.420 147.990 120.710 148.035 ;
        RECT 123.200 147.990 123.490 148.035 ;
        RECT 125.060 147.990 125.350 148.035 ;
        RECT 100.760 147.850 109.180 147.990 ;
        RECT 92.405 147.650 92.695 147.695 ;
        RECT 91.010 147.510 92.695 147.650 ;
        RECT 91.010 147.450 91.330 147.510 ;
        RECT 92.405 147.465 92.695 147.510 ;
        RECT 97.005 147.465 97.295 147.695 ;
        RECT 72.625 147.125 72.915 147.355 ;
        RECT 76.305 147.125 76.595 147.355 ;
        RECT 77.225 147.125 77.515 147.355 ;
        RECT 77.685 147.125 77.975 147.355 ;
        RECT 78.130 147.310 78.450 147.370 ;
        RECT 79.970 147.310 80.290 147.370 ;
        RECT 81.365 147.310 81.655 147.355 ;
        RECT 78.130 147.170 81.655 147.310 ;
        RECT 77.760 146.970 77.900 147.125 ;
        RECT 78.130 147.110 78.450 147.170 ;
        RECT 79.970 147.110 80.290 147.170 ;
        RECT 81.365 147.125 81.655 147.170 ;
        RECT 81.825 147.125 82.115 147.355 ;
        RECT 81.900 146.970 82.040 147.125 ;
        RECT 82.270 147.110 82.590 147.370 ;
        RECT 83.190 147.110 83.510 147.370 ;
        RECT 89.140 147.310 89.430 147.355 ;
        RECT 89.140 147.170 91.675 147.310 ;
        RECT 89.140 147.125 89.430 147.170 ;
        RECT 82.730 146.970 83.050 147.030 ;
        RECT 90.550 147.015 90.870 147.030 ;
        RECT 71.090 146.830 83.050 146.970 ;
        RECT 47.325 146.785 47.615 146.830 ;
        RECT 51.450 146.770 51.770 146.830 ;
        RECT 58.810 146.770 59.130 146.830 ;
        RECT 61.125 146.785 61.415 146.830 ;
        RECT 41.790 146.630 42.110 146.690 ;
        RECT 40.960 146.490 42.110 146.630 ;
        RECT 29.385 146.445 29.675 146.490 ;
        RECT 36.730 146.430 37.050 146.490 ;
        RECT 38.570 146.430 38.890 146.490 ;
        RECT 39.045 146.445 39.335 146.490 ;
        RECT 41.790 146.430 42.110 146.490 ;
        RECT 49.610 146.630 49.930 146.690 ;
        RECT 51.005 146.630 51.295 146.675 ;
        RECT 49.610 146.490 51.295 146.630 ;
        RECT 49.610 146.430 49.930 146.490 ;
        RECT 51.005 146.445 51.295 146.490 ;
        RECT 59.270 146.630 59.590 146.690 ;
        RECT 61.585 146.630 61.875 146.675 ;
        RECT 59.270 146.490 61.875 146.630 ;
        RECT 59.270 146.430 59.590 146.490 ;
        RECT 61.585 146.445 61.875 146.490 ;
        RECT 63.425 146.630 63.715 146.675 ;
        RECT 63.870 146.630 64.190 146.690 ;
        RECT 71.320 146.675 71.460 146.830 ;
        RECT 82.730 146.770 83.050 146.830 ;
        RECT 87.280 146.970 87.570 147.015 ;
        RECT 90.540 146.970 90.870 147.015 ;
        RECT 87.280 146.830 90.870 146.970 ;
        RECT 87.280 146.785 87.570 146.830 ;
        RECT 90.540 146.785 90.870 146.830 ;
        RECT 91.460 147.015 91.675 147.170 ;
        RECT 94.230 147.110 94.550 147.370 ;
        RECT 95.150 147.110 95.470 147.370 ;
        RECT 98.385 147.125 98.675 147.355 ;
        RECT 100.300 147.310 100.440 147.805 ;
        RECT 102.970 147.650 103.290 147.710 ;
        RECT 105.745 147.650 106.035 147.695 ;
        RECT 102.970 147.510 106.035 147.650 ;
        RECT 102.970 147.450 103.290 147.510 ;
        RECT 105.745 147.465 106.035 147.510 ;
        RECT 107.570 147.650 107.890 147.710 ;
        RECT 107.570 147.510 108.720 147.650 ;
        RECT 107.570 147.450 107.890 147.510 ;
        RECT 102.065 147.310 102.355 147.355 ;
        RECT 100.300 147.170 102.355 147.310 ;
        RECT 102.065 147.125 102.355 147.170 ;
        RECT 104.825 147.310 105.115 147.355 ;
        RECT 105.270 147.310 105.590 147.370 ;
        RECT 104.825 147.170 105.590 147.310 ;
        RECT 104.825 147.125 105.115 147.170 ;
        RECT 91.460 146.970 91.750 147.015 ;
        RECT 93.320 146.970 93.610 147.015 ;
        RECT 91.460 146.830 93.610 146.970 ;
        RECT 91.460 146.785 91.750 146.830 ;
        RECT 93.320 146.785 93.610 146.830 ;
        RECT 93.770 146.970 94.090 147.030 ;
        RECT 98.460 146.970 98.600 147.125 ;
        RECT 105.270 147.110 105.590 147.170 ;
        RECT 108.030 147.110 108.350 147.370 ;
        RECT 108.580 147.355 108.720 147.510 ;
        RECT 109.040 147.355 109.180 147.850 ;
        RECT 120.420 147.850 125.350 147.990 ;
        RECT 120.420 147.805 120.710 147.850 ;
        RECT 123.200 147.805 123.490 147.850 ;
        RECT 125.060 147.805 125.350 147.850 ;
        RECT 113.090 147.450 113.410 147.710 ;
        RECT 108.505 147.125 108.795 147.355 ;
        RECT 108.965 147.125 109.255 147.355 ;
        RECT 109.870 147.310 110.190 147.370 ;
        RECT 112.170 147.310 112.490 147.370 ;
        RECT 109.870 147.170 112.490 147.310 ;
        RECT 109.870 147.110 110.190 147.170 ;
        RECT 112.170 147.110 112.490 147.170 ;
        RECT 114.025 147.125 114.315 147.355 ;
        RECT 120.420 147.310 120.710 147.355 ;
        RECT 120.420 147.170 122.955 147.310 ;
        RECT 120.420 147.125 120.710 147.170 ;
        RECT 93.770 146.830 98.600 146.970 ;
        RECT 106.205 146.970 106.495 147.015 ;
        RECT 106.665 146.970 106.955 147.015 ;
        RECT 114.100 146.970 114.240 147.125 ;
        RECT 106.205 146.830 106.955 146.970 ;
        RECT 90.550 146.770 90.870 146.785 ;
        RECT 93.770 146.770 94.090 146.830 ;
        RECT 106.205 146.785 106.495 146.830 ;
        RECT 106.665 146.785 106.955 146.830 ;
        RECT 107.200 146.830 114.240 146.970 ;
        RECT 116.555 146.970 116.845 147.015 ;
        RECT 117.690 146.970 118.010 147.030 ;
        RECT 116.555 146.830 118.010 146.970 ;
        RECT 63.425 146.490 64.190 146.630 ;
        RECT 63.425 146.445 63.715 146.490 ;
        RECT 63.870 146.430 64.190 146.490 ;
        RECT 71.245 146.445 71.535 146.675 ;
        RECT 73.530 146.630 73.850 146.690 ;
        RECT 78.130 146.630 78.450 146.690 ;
        RECT 73.530 146.490 78.450 146.630 ;
        RECT 73.530 146.430 73.850 146.490 ;
        RECT 78.130 146.430 78.450 146.490 ;
        RECT 79.510 146.430 79.830 146.690 ;
        RECT 82.270 146.630 82.590 146.690 ;
        RECT 85.275 146.630 85.565 146.675 ;
        RECT 85.950 146.630 86.270 146.690 ;
        RECT 82.270 146.490 86.270 146.630 ;
        RECT 82.270 146.430 82.590 146.490 ;
        RECT 85.275 146.445 85.565 146.490 ;
        RECT 85.950 146.430 86.270 146.490 ;
        RECT 96.990 146.630 97.310 146.690 ;
        RECT 97.925 146.630 98.215 146.675 ;
        RECT 107.200 146.630 107.340 146.830 ;
        RECT 116.555 146.785 116.845 146.830 ;
        RECT 117.690 146.770 118.010 146.830 ;
        RECT 118.560 146.970 118.850 147.015 ;
        RECT 119.990 146.970 120.310 147.030 ;
        RECT 122.740 147.015 122.955 147.170 ;
        RECT 123.670 147.110 123.990 147.370 ;
        RECT 125.525 147.310 125.815 147.355 ;
        RECT 125.970 147.310 126.290 147.370 ;
        RECT 125.525 147.170 126.290 147.310 ;
        RECT 125.525 147.125 125.815 147.170 ;
        RECT 125.970 147.110 126.290 147.170 ;
        RECT 121.820 146.970 122.110 147.015 ;
        RECT 118.560 146.830 122.110 146.970 ;
        RECT 118.560 146.785 118.850 146.830 ;
        RECT 119.990 146.770 120.310 146.830 ;
        RECT 121.820 146.785 122.110 146.830 ;
        RECT 122.740 146.970 123.030 147.015 ;
        RECT 124.600 146.970 124.890 147.015 ;
        RECT 122.740 146.830 124.890 146.970 ;
        RECT 122.740 146.785 123.030 146.830 ;
        RECT 124.600 146.785 124.890 146.830 ;
        RECT 96.990 146.490 107.340 146.630 ;
        RECT 108.030 146.630 108.350 146.690 ;
        RECT 109.410 146.630 109.730 146.690 ;
        RECT 108.030 146.490 109.730 146.630 ;
        RECT 96.990 146.430 97.310 146.490 ;
        RECT 97.925 146.445 98.215 146.490 ;
        RECT 108.030 146.430 108.350 146.490 ;
        RECT 109.410 146.430 109.730 146.490 ;
        RECT 113.565 146.630 113.855 146.675 ;
        RECT 114.010 146.630 114.330 146.690 ;
        RECT 117.230 146.630 117.550 146.690 ;
        RECT 113.565 146.490 117.550 146.630 ;
        RECT 113.565 146.445 113.855 146.490 ;
        RECT 114.010 146.430 114.330 146.490 ;
        RECT 117.230 146.430 117.550 146.490 ;
        RECT 14.580 145.810 127.740 146.290 ;
        RECT 20.170 145.410 20.490 145.670 ;
        RECT 22.930 145.655 23.250 145.670 ;
        RECT 22.715 145.425 23.250 145.655 ;
        RECT 50.990 145.610 51.310 145.670 ;
        RECT 22.930 145.410 23.250 145.425 ;
        RECT 40.960 145.470 51.310 145.610 ;
        RECT 21.565 145.270 21.855 145.315 ;
        RECT 24.720 145.270 25.010 145.315 ;
        RECT 27.980 145.270 28.270 145.315 ;
        RECT 21.565 145.130 28.270 145.270 ;
        RECT 21.565 145.085 21.855 145.130 ;
        RECT 24.720 145.085 25.010 145.130 ;
        RECT 27.980 145.085 28.270 145.130 ;
        RECT 28.900 145.270 29.190 145.315 ;
        RECT 30.760 145.270 31.050 145.315 ;
        RECT 28.900 145.130 31.050 145.270 ;
        RECT 28.900 145.085 29.190 145.130 ;
        RECT 30.760 145.085 31.050 145.130 ;
        RECT 19.725 144.930 20.015 144.975 ;
        RECT 21.105 144.930 21.395 144.975 ;
        RECT 19.725 144.790 21.395 144.930 ;
        RECT 19.725 144.745 20.015 144.790 ;
        RECT 21.105 144.745 21.395 144.790 ;
        RECT 26.580 144.930 26.870 144.975 ;
        RECT 28.900 144.930 29.115 145.085 ;
        RECT 26.580 144.790 29.115 144.930 ;
        RECT 30.290 144.930 30.610 144.990 ;
        RECT 40.960 144.975 41.100 145.470 ;
        RECT 50.990 145.410 51.310 145.470 ;
        RECT 51.910 145.410 52.230 145.670 ;
        RECT 53.750 145.410 54.070 145.670 ;
        RECT 80.890 145.610 81.210 145.670 ;
        RECT 80.520 145.470 81.210 145.610 ;
        RECT 41.345 145.270 41.635 145.315 ;
        RECT 44.500 145.270 44.790 145.315 ;
        RECT 47.760 145.270 48.050 145.315 ;
        RECT 41.345 145.130 48.050 145.270 ;
        RECT 41.345 145.085 41.635 145.130 ;
        RECT 44.500 145.085 44.790 145.130 ;
        RECT 47.760 145.085 48.050 145.130 ;
        RECT 48.680 145.270 48.970 145.315 ;
        RECT 50.540 145.270 50.830 145.315 ;
        RECT 48.680 145.130 50.830 145.270 ;
        RECT 51.080 145.270 51.220 145.410 ;
        RECT 55.130 145.270 55.450 145.330 ;
        RECT 59.270 145.270 59.590 145.330 ;
        RECT 65.265 145.270 65.555 145.315 ;
        RECT 51.080 145.130 58.580 145.270 ;
        RECT 48.680 145.085 48.970 145.130 ;
        RECT 50.540 145.085 50.830 145.130 ;
        RECT 40.885 144.930 41.175 144.975 ;
        RECT 30.290 144.790 41.175 144.930 ;
        RECT 26.580 144.745 26.870 144.790 ;
        RECT 21.180 143.910 21.320 144.745 ;
        RECT 30.290 144.730 30.610 144.790 ;
        RECT 40.885 144.745 41.175 144.790 ;
        RECT 46.360 144.930 46.650 144.975 ;
        RECT 48.680 144.930 48.895 145.085 ;
        RECT 55.130 145.070 55.450 145.130 ;
        RECT 46.360 144.790 48.895 144.930 ;
        RECT 46.360 144.745 46.650 144.790 ;
        RECT 49.610 144.730 49.930 144.990 ;
        RECT 58.440 144.975 58.580 145.130 ;
        RECT 59.270 145.130 65.555 145.270 ;
        RECT 59.270 145.070 59.590 145.130 ;
        RECT 65.265 145.085 65.555 145.130 ;
        RECT 79.510 145.070 79.830 145.330 ;
        RECT 54.225 144.930 54.515 144.975 ;
        RECT 50.160 144.790 54.515 144.930 ;
        RECT 28.910 144.590 29.230 144.650 ;
        RECT 29.845 144.590 30.135 144.635 ;
        RECT 28.910 144.450 30.135 144.590 ;
        RECT 28.910 144.390 29.230 144.450 ;
        RECT 29.845 144.405 30.135 144.450 ;
        RECT 31.685 144.590 31.975 144.635 ;
        RECT 36.270 144.590 36.590 144.650 ;
        RECT 31.685 144.450 36.590 144.590 ;
        RECT 31.685 144.405 31.975 144.450 ;
        RECT 36.270 144.390 36.590 144.450 ;
        RECT 42.495 144.590 42.785 144.635 ;
        RECT 50.160 144.590 50.300 144.790 ;
        RECT 54.225 144.745 54.515 144.790 ;
        RECT 58.365 144.745 58.655 144.975 ;
        RECT 65.710 144.730 66.030 144.990 ;
        RECT 80.520 144.975 80.660 145.470 ;
        RECT 80.890 145.410 81.210 145.470 ;
        RECT 85.950 145.410 86.270 145.670 ;
        RECT 91.010 145.410 91.330 145.670 ;
        RECT 96.990 145.410 97.310 145.670 ;
        RECT 117.230 145.410 117.550 145.670 ;
        RECT 119.990 145.410 120.310 145.670 ;
        RECT 122.305 145.610 122.595 145.655 ;
        RECT 123.670 145.610 123.990 145.670 ;
        RECT 122.305 145.470 123.990 145.610 ;
        RECT 122.305 145.425 122.595 145.470 ;
        RECT 123.670 145.410 123.990 145.470 ;
        RECT 107.125 145.270 107.415 145.315 ;
        RECT 109.885 145.270 110.175 145.315 ;
        RECT 107.125 145.130 110.175 145.270 ;
        RECT 107.125 145.085 107.415 145.130 ;
        RECT 109.885 145.085 110.175 145.130 ;
        RECT 112.260 145.130 117.000 145.270 ;
        RECT 80.445 144.745 80.735 144.975 ;
        RECT 80.905 144.930 81.195 144.975 ;
        RECT 81.350 144.930 81.670 144.990 ;
        RECT 80.905 144.790 81.670 144.930 ;
        RECT 80.905 144.745 81.195 144.790 ;
        RECT 81.350 144.730 81.670 144.790 ;
        RECT 84.570 144.930 84.890 144.990 ;
        RECT 86.425 144.930 86.715 144.975 ;
        RECT 90.105 144.930 90.395 144.975 ;
        RECT 84.570 144.790 86.715 144.930 ;
        RECT 84.570 144.730 84.890 144.790 ;
        RECT 86.425 144.745 86.715 144.790 ;
        RECT 88.340 144.790 90.395 144.930 ;
        RECT 50.530 144.590 50.850 144.650 ;
        RECT 42.495 144.450 50.850 144.590 ;
        RECT 42.495 144.405 42.785 144.450 ;
        RECT 50.530 144.390 50.850 144.450 ;
        RECT 51.465 144.405 51.755 144.635 ;
        RECT 54.670 144.590 54.990 144.650 ;
        RECT 55.145 144.590 55.435 144.635 ;
        RECT 64.790 144.590 65.110 144.650 ;
        RECT 69.390 144.590 69.710 144.650 ;
        RECT 54.670 144.450 69.710 144.590 ;
        RECT 26.580 144.250 26.870 144.295 ;
        RECT 29.360 144.250 29.650 144.295 ;
        RECT 31.220 144.250 31.510 144.295 ;
        RECT 26.580 144.110 31.510 144.250 ;
        RECT 26.580 144.065 26.870 144.110 ;
        RECT 29.360 144.065 29.650 144.110 ;
        RECT 31.220 144.065 31.510 144.110 ;
        RECT 46.360 144.250 46.650 144.295 ;
        RECT 49.140 144.250 49.430 144.295 ;
        RECT 51.000 144.250 51.290 144.295 ;
        RECT 46.360 144.110 51.290 144.250 ;
        RECT 51.540 144.250 51.680 144.405 ;
        RECT 54.670 144.390 54.990 144.450 ;
        RECT 55.145 144.405 55.435 144.450 ;
        RECT 64.790 144.390 65.110 144.450 ;
        RECT 69.390 144.390 69.710 144.450 ;
        RECT 85.030 144.390 85.350 144.650 ;
        RECT 63.870 144.250 64.190 144.310 ;
        RECT 51.540 144.110 64.190 144.250 ;
        RECT 46.360 144.065 46.650 144.110 ;
        RECT 49.140 144.065 49.430 144.110 ;
        RECT 51.000 144.065 51.290 144.110 ;
        RECT 63.870 144.050 64.190 144.110 ;
        RECT 68.930 144.250 69.250 144.310 ;
        RECT 70.770 144.250 71.090 144.310 ;
        RECT 68.930 144.110 71.090 144.250 ;
        RECT 68.930 144.050 69.250 144.110 ;
        RECT 70.770 144.050 71.090 144.110 ;
        RECT 75.370 144.250 75.690 144.310 ;
        RECT 88.340 144.295 88.480 144.790 ;
        RECT 90.105 144.745 90.395 144.790 ;
        RECT 94.245 144.930 94.535 144.975 ;
        RECT 96.530 144.930 96.850 144.990 ;
        RECT 94.245 144.790 96.850 144.930 ;
        RECT 94.245 144.745 94.535 144.790 ;
        RECT 96.530 144.730 96.850 144.790 ;
        RECT 108.505 144.930 108.795 144.975 ;
        RECT 108.950 144.930 109.270 144.990 ;
        RECT 108.505 144.790 109.270 144.930 ;
        RECT 108.505 144.745 108.795 144.790 ;
        RECT 108.950 144.730 109.270 144.790 ;
        RECT 109.410 144.930 109.730 144.990 ;
        RECT 111.265 144.930 111.555 144.975 ;
        RECT 109.410 144.790 111.555 144.930 ;
        RECT 109.410 144.730 109.730 144.790 ;
        RECT 111.265 144.745 111.555 144.790 ;
        RECT 108.045 144.590 108.335 144.635 ;
        RECT 110.330 144.590 110.650 144.650 ;
        RECT 108.045 144.450 110.650 144.590 ;
        RECT 108.045 144.405 108.335 144.450 ;
        RECT 110.330 144.390 110.650 144.450 ;
        RECT 81.825 144.250 82.115 144.295 ;
        RECT 75.370 144.110 82.115 144.250 ;
        RECT 75.370 144.050 75.690 144.110 ;
        RECT 81.825 144.065 82.115 144.110 ;
        RECT 88.265 144.065 88.555 144.295 ;
        RECT 108.950 144.250 109.270 144.310 ;
        RECT 109.425 144.250 109.715 144.295 ;
        RECT 111.340 144.250 111.480 144.745 ;
        RECT 111.710 144.730 112.030 144.990 ;
        RECT 112.260 144.975 112.400 145.130 ;
        RECT 112.185 144.745 112.475 144.975 ;
        RECT 112.630 144.930 112.950 144.990 ;
        RECT 113.105 144.930 113.395 144.975 ;
        RECT 112.630 144.790 113.395 144.930 ;
        RECT 112.630 144.730 112.950 144.790 ;
        RECT 113.105 144.745 113.395 144.790 ;
        RECT 113.550 144.590 113.870 144.650 ;
        RECT 116.860 144.635 117.000 145.130 ;
        RECT 119.530 144.730 119.850 144.990 ;
        RECT 121.385 144.745 121.675 144.975 ;
        RECT 115.865 144.590 116.155 144.635 ;
        RECT 113.550 144.450 116.155 144.590 ;
        RECT 113.550 144.390 113.870 144.450 ;
        RECT 115.865 144.405 116.155 144.450 ;
        RECT 116.785 144.590 117.075 144.635 ;
        RECT 117.690 144.590 118.010 144.650 ;
        RECT 121.460 144.590 121.600 144.745 ;
        RECT 116.785 144.450 118.010 144.590 ;
        RECT 116.785 144.405 117.075 144.450 ;
        RECT 117.690 144.390 118.010 144.450 ;
        RECT 119.160 144.450 121.600 144.590 ;
        RECT 119.160 144.295 119.300 144.450 ;
        RECT 108.950 144.110 109.715 144.250 ;
        RECT 108.950 144.050 109.270 144.110 ;
        RECT 109.425 144.065 109.715 144.110 ;
        RECT 110.420 144.110 111.480 144.250 ;
        RECT 110.420 143.970 110.560 144.110 ;
        RECT 119.085 144.065 119.375 144.295 ;
        RECT 29.830 143.910 30.150 143.970 ;
        RECT 21.180 143.770 30.150 143.910 ;
        RECT 29.830 143.710 30.150 143.770 ;
        RECT 58.810 143.710 59.130 143.970 ;
        RECT 67.565 143.910 67.855 143.955 ;
        RECT 69.850 143.910 70.170 143.970 ;
        RECT 67.565 143.770 70.170 143.910 ;
        RECT 67.565 143.725 67.855 143.770 ;
        RECT 69.850 143.710 70.170 143.770 ;
        RECT 80.890 143.710 81.210 143.970 ;
        RECT 108.505 143.910 108.795 143.955 ;
        RECT 109.870 143.910 110.190 143.970 ;
        RECT 108.505 143.770 110.190 143.910 ;
        RECT 108.505 143.725 108.795 143.770 ;
        RECT 109.870 143.710 110.190 143.770 ;
        RECT 110.330 143.710 110.650 143.970 ;
        RECT 14.580 143.090 127.740 143.570 ;
        RECT 35.810 142.690 36.130 142.950 ;
        RECT 48.245 142.705 48.535 142.935 ;
        RECT 45.010 142.550 45.330 142.610 ;
        RECT 48.320 142.550 48.460 142.705 ;
        RECT 59.270 142.690 59.590 142.950 ;
        RECT 108.950 142.890 109.270 142.950 ;
        RECT 111.710 142.890 112.030 142.950 ;
        RECT 108.950 142.750 112.030 142.890 ;
        RECT 108.950 142.690 109.270 142.750 ;
        RECT 111.710 142.690 112.030 142.750 ;
        RECT 45.010 142.410 48.460 142.550 ;
        RECT 62.605 142.550 62.895 142.595 ;
        RECT 65.725 142.550 66.015 142.595 ;
        RECT 67.615 142.550 67.905 142.595 ;
        RECT 68.930 142.550 69.250 142.610 ;
        RECT 62.605 142.410 67.905 142.550 ;
        RECT 45.010 142.350 45.330 142.410 ;
        RECT 62.605 142.365 62.895 142.410 ;
        RECT 65.725 142.365 66.015 142.410 ;
        RECT 67.615 142.365 67.905 142.410 ;
        RECT 68.100 142.410 69.250 142.550 ;
        RECT 34.430 142.210 34.750 142.270 ;
        RECT 35.825 142.210 36.115 142.255 ;
        RECT 34.430 142.070 36.115 142.210 ;
        RECT 34.430 142.010 34.750 142.070 ;
        RECT 35.825 142.025 36.115 142.070 ;
        RECT 46.390 142.210 46.710 142.270 ;
        RECT 48.705 142.210 48.995 142.255 ;
        RECT 46.390 142.070 48.995 142.210 ;
        RECT 46.390 142.010 46.710 142.070 ;
        RECT 48.705 142.025 48.995 142.070 ;
        RECT 53.290 142.210 53.610 142.270 ;
        RECT 56.525 142.210 56.815 142.255 ;
        RECT 59.745 142.210 60.035 142.255 ;
        RECT 68.100 142.210 68.240 142.410 ;
        RECT 68.930 142.350 69.250 142.410 ;
        RECT 53.290 142.070 54.440 142.210 ;
        RECT 53.290 142.010 53.610 142.070 ;
        RECT 34.890 141.870 35.210 141.930 ;
        RECT 35.365 141.870 35.655 141.915 ;
        RECT 34.890 141.730 35.655 141.870 ;
        RECT 34.890 141.670 35.210 141.730 ;
        RECT 35.365 141.685 35.655 141.730 ;
        RECT 45.930 141.870 46.250 141.930 ;
        RECT 48.245 141.870 48.535 141.915 ;
        RECT 45.930 141.730 48.535 141.870 ;
        RECT 45.930 141.670 46.250 141.730 ;
        RECT 48.245 141.685 48.535 141.730 ;
        RECT 53.750 141.670 54.070 141.930 ;
        RECT 54.300 141.915 54.440 142.070 ;
        RECT 54.760 142.070 60.035 142.210 ;
        RECT 54.760 141.915 54.900 142.070 ;
        RECT 56.525 142.025 56.815 142.070 ;
        RECT 59.745 142.025 60.035 142.070 ;
        RECT 60.280 142.070 68.240 142.210 ;
        RECT 54.225 141.685 54.515 141.915 ;
        RECT 54.685 141.685 54.975 141.915 ;
        RECT 55.605 141.870 55.895 141.915 ;
        RECT 56.050 141.870 56.370 141.930 ;
        RECT 60.280 141.870 60.420 142.070 ;
        RECT 68.470 142.010 68.790 142.270 ;
        RECT 113.090 142.210 113.410 142.270 ;
        RECT 116.325 142.210 116.615 142.255 ;
        RECT 113.090 142.070 116.615 142.210 ;
        RECT 113.090 142.010 113.410 142.070 ;
        RECT 116.325 142.025 116.615 142.070 ;
        RECT 55.605 141.730 56.370 141.870 ;
        RECT 55.605 141.685 55.895 141.730 ;
        RECT 56.050 141.670 56.370 141.730 ;
        RECT 57.980 141.730 60.420 141.870 ;
        RECT 36.745 141.530 37.035 141.575 ;
        RECT 39.490 141.530 39.810 141.590 ;
        RECT 36.745 141.390 39.810 141.530 ;
        RECT 36.745 141.345 37.035 141.390 ;
        RECT 39.490 141.330 39.810 141.390 ;
        RECT 49.625 141.530 49.915 141.575 ;
        RECT 52.385 141.530 52.675 141.575 ;
        RECT 49.625 141.390 52.675 141.530 ;
        RECT 49.625 141.345 49.915 141.390 ;
        RECT 52.385 141.345 52.675 141.390 ;
        RECT 29.370 141.190 29.690 141.250 ;
        RECT 34.445 141.190 34.735 141.235 ;
        RECT 29.370 141.050 34.735 141.190 ;
        RECT 29.370 140.990 29.690 141.050 ;
        RECT 34.445 141.005 34.735 141.050 ;
        RECT 47.325 141.190 47.615 141.235 ;
        RECT 57.980 141.190 58.120 141.730 ;
        RECT 58.810 141.530 59.130 141.590 ;
        RECT 61.525 141.575 61.815 141.890 ;
        RECT 62.605 141.870 62.895 141.915 ;
        RECT 66.185 141.870 66.475 141.915 ;
        RECT 68.020 141.870 68.310 141.915 ;
        RECT 62.605 141.730 68.310 141.870 ;
        RECT 62.605 141.685 62.895 141.730 ;
        RECT 66.185 141.685 66.475 141.730 ;
        RECT 68.020 141.685 68.310 141.730 ;
        RECT 69.850 141.670 70.170 141.930 ;
        RECT 70.770 141.870 71.090 141.930 ;
        RECT 72.625 141.870 72.915 141.915 ;
        RECT 70.770 141.730 72.915 141.870 ;
        RECT 70.770 141.670 71.090 141.730 ;
        RECT 72.625 141.685 72.915 141.730 ;
        RECT 117.690 141.670 118.010 141.930 ;
        RECT 119.530 141.870 119.850 141.930 ;
        RECT 120.005 141.870 120.295 141.915 ;
        RECT 119.530 141.730 120.295 141.870 ;
        RECT 119.530 141.670 119.850 141.730 ;
        RECT 120.005 141.685 120.295 141.730 ;
        RECT 61.225 141.530 61.815 141.575 ;
        RECT 64.465 141.530 65.115 141.575 ;
        RECT 58.810 141.390 65.115 141.530 ;
        RECT 58.810 141.330 59.130 141.390 ;
        RECT 61.225 141.345 61.515 141.390 ;
        RECT 64.465 141.345 65.115 141.390 ;
        RECT 67.105 141.530 67.395 141.575 ;
        RECT 67.105 141.390 69.160 141.530 ;
        RECT 67.105 141.345 67.395 141.390 ;
        RECT 47.325 141.050 58.120 141.190 ;
        RECT 63.870 141.190 64.190 141.250 ;
        RECT 68.470 141.190 68.790 141.250 ;
        RECT 69.020 141.235 69.160 141.390 ;
        RECT 63.870 141.050 68.790 141.190 ;
        RECT 47.325 141.005 47.615 141.050 ;
        RECT 63.870 140.990 64.190 141.050 ;
        RECT 68.470 140.990 68.790 141.050 ;
        RECT 68.945 141.005 69.235 141.235 ;
        RECT 72.150 140.990 72.470 141.250 ;
        RECT 117.230 140.990 117.550 141.250 ;
        RECT 119.530 140.990 119.850 141.250 ;
        RECT 120.450 140.990 120.770 141.250 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 14.580 140.370 127.740 140.850 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 35.810 139.970 36.130 140.230 ;
        RECT 38.585 139.985 38.875 140.215 ;
        RECT 39.490 140.170 39.810 140.230 ;
        RECT 59.285 140.170 59.575 140.215 ;
        RECT 61.110 140.170 61.430 140.230 ;
        RECT 63.885 140.170 64.175 140.215 ;
        RECT 39.490 140.030 59.575 140.170 ;
        RECT 18.280 139.830 18.570 139.875 ;
        RECT 19.250 139.830 19.570 139.890 ;
        RECT 21.540 139.830 21.830 139.875 ;
        RECT 18.280 139.690 21.830 139.830 ;
        RECT 18.280 139.645 18.570 139.690 ;
        RECT 19.250 139.630 19.570 139.690 ;
        RECT 21.540 139.645 21.830 139.690 ;
        RECT 22.460 139.830 22.750 139.875 ;
        RECT 24.320 139.830 24.610 139.875 ;
        RECT 38.660 139.830 38.800 139.985 ;
        RECT 39.490 139.970 39.810 140.030 ;
        RECT 59.285 139.985 59.575 140.030 ;
        RECT 59.820 140.030 64.175 140.170 ;
        RECT 22.460 139.690 24.610 139.830 ;
        RECT 22.460 139.645 22.750 139.690 ;
        RECT 24.320 139.645 24.610 139.690 ;
        RECT 36.590 139.690 38.800 139.830 ;
        RECT 40.885 139.830 41.175 139.875 ;
        RECT 41.330 139.830 41.650 139.890 ;
        RECT 59.820 139.830 59.960 140.030 ;
        RECT 61.110 139.970 61.430 140.030 ;
        RECT 63.885 139.985 64.175 140.030 ;
        RECT 65.710 140.170 66.030 140.230 ;
        RECT 67.795 140.170 68.085 140.215 ;
        RECT 65.710 140.030 68.085 140.170 ;
        RECT 65.710 139.970 66.030 140.030 ;
        RECT 67.795 139.985 68.085 140.030 ;
        RECT 81.350 139.970 81.670 140.230 ;
        RECT 84.570 140.170 84.890 140.230 ;
        RECT 85.965 140.170 86.255 140.215 ;
        RECT 84.570 140.030 86.255 140.170 ;
        RECT 84.570 139.970 84.890 140.030 ;
        RECT 85.965 139.985 86.255 140.030 ;
        RECT 88.265 139.985 88.555 140.215 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 65.800 139.830 65.940 139.970 ;
        RECT 40.885 139.690 41.650 139.830 ;
        RECT 20.140 139.490 20.430 139.535 ;
        RECT 22.460 139.490 22.675 139.645 ;
        RECT 20.140 139.350 22.675 139.490 ;
        RECT 34.890 139.490 35.210 139.550 ;
        RECT 35.810 139.490 36.130 139.550 ;
        RECT 36.590 139.490 36.730 139.690 ;
        RECT 40.885 139.645 41.175 139.690 ;
        RECT 41.330 139.630 41.650 139.690 ;
        RECT 55.220 139.690 59.960 139.830 ;
        RECT 61.660 139.690 65.940 139.830 ;
        RECT 69.800 139.830 70.090 139.875 ;
        RECT 72.150 139.830 72.470 139.890 ;
        RECT 73.060 139.830 73.350 139.875 ;
        RECT 69.800 139.690 73.350 139.830 ;
        RECT 34.890 139.350 35.405 139.490 ;
        RECT 35.810 139.350 36.730 139.490 ;
        RECT 39.505 139.490 39.795 139.535 ;
        RECT 55.220 139.490 55.360 139.690 ;
        RECT 39.505 139.350 55.360 139.490 ;
        RECT 20.140 139.305 20.430 139.350 ;
        RECT 34.890 139.290 35.210 139.350 ;
        RECT 35.810 139.290 36.130 139.350 ;
        RECT 39.505 139.305 39.795 139.350 ;
        RECT 55.605 139.305 55.895 139.535 ;
        RECT 23.390 138.950 23.710 139.210 ;
        RECT 25.245 139.150 25.535 139.195 ;
        RECT 29.830 139.150 30.150 139.210 ;
        RECT 25.245 139.010 30.150 139.150 ;
        RECT 25.245 138.965 25.535 139.010 ;
        RECT 29.830 138.950 30.150 139.010 ;
        RECT 30.290 139.150 30.610 139.210 ;
        RECT 33.985 139.150 34.275 139.195 ;
        RECT 30.290 139.010 34.275 139.150 ;
        RECT 30.290 138.950 30.610 139.010 ;
        RECT 33.985 138.965 34.275 139.010 ;
        RECT 39.950 138.950 40.270 139.210 ;
        RECT 55.130 139.150 55.450 139.210 ;
        RECT 55.680 139.150 55.820 139.305 ;
        RECT 56.050 139.290 56.370 139.550 ;
        RECT 60.650 139.290 60.970 139.550 ;
        RECT 61.660 139.535 61.800 139.690 ;
        RECT 69.800 139.645 70.090 139.690 ;
        RECT 72.150 139.630 72.470 139.690 ;
        RECT 73.060 139.645 73.350 139.690 ;
        RECT 73.980 139.830 74.270 139.875 ;
        RECT 75.840 139.830 76.130 139.875 ;
        RECT 73.980 139.690 76.130 139.830 ;
        RECT 73.980 139.645 74.270 139.690 ;
        RECT 75.840 139.645 76.130 139.690 ;
        RECT 79.970 139.830 80.290 139.890 ;
        RECT 81.440 139.830 81.580 139.970 ;
        RECT 84.660 139.830 84.800 139.970 ;
        RECT 79.970 139.690 81.580 139.830 ;
        RECT 81.900 139.690 84.800 139.830 ;
        RECT 61.125 139.305 61.415 139.535 ;
        RECT 61.585 139.305 61.875 139.535 ;
        RECT 62.505 139.305 62.795 139.535 ;
        RECT 55.130 139.010 55.820 139.150 ;
        RECT 55.130 138.950 55.450 139.010 ;
        RECT 20.140 138.810 20.430 138.855 ;
        RECT 22.920 138.810 23.210 138.855 ;
        RECT 24.780 138.810 25.070 138.855 ;
        RECT 20.140 138.670 25.070 138.810 ;
        RECT 20.140 138.625 20.430 138.670 ;
        RECT 22.920 138.625 23.210 138.670 ;
        RECT 24.780 138.625 25.070 138.670 ;
        RECT 16.275 138.470 16.565 138.515 ;
        RECT 22.470 138.470 22.790 138.530 ;
        RECT 16.275 138.330 22.790 138.470 ;
        RECT 16.275 138.285 16.565 138.330 ;
        RECT 22.470 138.270 22.790 138.330 ;
        RECT 34.430 138.470 34.750 138.530 ;
        RECT 39.505 138.470 39.795 138.515 ;
        RECT 34.430 138.330 39.795 138.470 ;
        RECT 34.430 138.270 34.750 138.330 ;
        RECT 39.505 138.285 39.795 138.330 ;
        RECT 47.770 138.470 48.090 138.530 ;
        RECT 50.070 138.470 50.390 138.530 ;
        RECT 53.750 138.470 54.070 138.530 ;
        RECT 47.770 138.330 54.070 138.470 ;
        RECT 61.200 138.470 61.340 139.305 ;
        RECT 62.580 138.810 62.720 139.305 ;
        RECT 65.250 139.290 65.570 139.550 ;
        RECT 65.725 139.305 66.015 139.535 ;
        RECT 65.800 139.150 65.940 139.305 ;
        RECT 66.170 139.290 66.490 139.550 ;
        RECT 67.105 139.490 67.395 139.535 ;
        RECT 68.010 139.490 68.330 139.550 ;
        RECT 67.105 139.350 68.330 139.490 ;
        RECT 67.105 139.305 67.395 139.350 ;
        RECT 68.010 139.290 68.330 139.350 ;
        RECT 71.660 139.490 71.950 139.535 ;
        RECT 73.980 139.490 74.195 139.645 ;
        RECT 79.970 139.630 80.290 139.690 ;
        RECT 80.980 139.535 81.120 139.690 ;
        RECT 81.900 139.535 82.040 139.690 ;
        RECT 71.660 139.350 74.195 139.490 ;
        RECT 71.660 139.305 71.950 139.350 ;
        RECT 80.905 139.305 81.195 139.535 ;
        RECT 81.365 139.305 81.655 139.535 ;
        RECT 81.825 139.305 82.115 139.535 ;
        RECT 82.745 139.305 83.035 139.535 ;
        RECT 70.310 139.150 70.630 139.210 ;
        RECT 65.800 139.010 70.630 139.150 ;
        RECT 64.330 138.810 64.650 138.870 ;
        RECT 67.550 138.810 67.870 138.870 ;
        RECT 62.580 138.670 67.870 138.810 ;
        RECT 64.330 138.610 64.650 138.670 ;
        RECT 67.550 138.610 67.870 138.670 ;
        RECT 66.630 138.470 66.950 138.530 ;
        RECT 68.100 138.470 68.240 139.010 ;
        RECT 70.310 138.950 70.630 139.010 ;
        RECT 74.910 138.950 75.230 139.210 ;
        RECT 76.765 138.965 77.055 139.195 ;
        RECT 81.440 139.150 81.580 139.305 ;
        RECT 82.270 139.150 82.590 139.210 ;
        RECT 81.440 139.010 82.590 139.150 ;
        RECT 82.820 139.150 82.960 139.305 ;
        RECT 86.410 139.290 86.730 139.550 ;
        RECT 88.340 139.490 88.480 139.985 ;
        RECT 100.160 139.830 100.450 139.875 ;
        RECT 102.510 139.830 102.830 139.890 ;
        RECT 103.420 139.830 103.710 139.875 ;
        RECT 100.160 139.690 103.710 139.830 ;
        RECT 100.160 139.645 100.450 139.690 ;
        RECT 102.510 139.630 102.830 139.690 ;
        RECT 103.420 139.645 103.710 139.690 ;
        RECT 104.340 139.830 104.630 139.875 ;
        RECT 106.200 139.830 106.490 139.875 ;
        RECT 104.340 139.690 106.490 139.830 ;
        RECT 104.340 139.645 104.630 139.690 ;
        RECT 106.200 139.645 106.490 139.690 ;
        RECT 110.330 139.830 110.650 139.890 ;
        RECT 112.170 139.830 112.490 139.890 ;
        RECT 117.230 139.875 117.550 139.890 ;
        RECT 113.105 139.830 113.395 139.875 ;
        RECT 117.015 139.830 117.550 139.875 ;
        RECT 110.330 139.690 111.940 139.830 ;
        RECT 89.185 139.490 89.475 139.535 ;
        RECT 88.340 139.350 89.475 139.490 ;
        RECT 89.185 139.305 89.475 139.350 ;
        RECT 102.020 139.490 102.310 139.535 ;
        RECT 104.340 139.490 104.555 139.645 ;
        RECT 110.330 139.630 110.650 139.690 ;
        RECT 102.020 139.350 104.555 139.490 ;
        RECT 109.410 139.490 109.730 139.550 ;
        RECT 109.885 139.490 110.175 139.535 ;
        RECT 109.410 139.350 110.175 139.490 ;
        RECT 110.805 139.480 111.095 139.550 ;
        RECT 111.800 139.535 111.940 139.690 ;
        RECT 112.170 139.690 113.395 139.830 ;
        RECT 112.170 139.630 112.490 139.690 ;
        RECT 113.105 139.645 113.395 139.690 ;
        RECT 114.100 139.690 117.550 139.830 ;
        RECT 102.020 139.305 102.310 139.350 ;
        RECT 109.410 139.290 109.730 139.350 ;
        RECT 109.885 139.305 110.175 139.350 ;
        RECT 110.420 139.340 111.095 139.480 ;
        RECT 83.190 139.150 83.510 139.210 ;
        RECT 82.820 139.010 83.510 139.150 ;
        RECT 71.660 138.810 71.950 138.855 ;
        RECT 74.440 138.810 74.730 138.855 ;
        RECT 76.300 138.810 76.590 138.855 ;
        RECT 71.660 138.670 76.590 138.810 ;
        RECT 76.840 138.810 76.980 138.965 ;
        RECT 82.270 138.950 82.590 139.010 ;
        RECT 83.190 138.950 83.510 139.010 ;
        RECT 85.030 138.950 85.350 139.210 ;
        RECT 98.155 139.150 98.445 139.195 ;
        RECT 98.830 139.150 99.150 139.210 ;
        RECT 98.155 139.010 99.150 139.150 ;
        RECT 98.155 138.965 98.445 139.010 ;
        RECT 98.830 138.950 99.150 139.010 ;
        RECT 105.270 138.950 105.590 139.210 ;
        RECT 107.125 138.965 107.415 139.195 ;
        RECT 94.230 138.810 94.550 138.870 ;
        RECT 76.840 138.670 94.550 138.810 ;
        RECT 71.660 138.625 71.950 138.670 ;
        RECT 74.440 138.625 74.730 138.670 ;
        RECT 76.300 138.625 76.590 138.670 ;
        RECT 94.230 138.610 94.550 138.670 ;
        RECT 102.020 138.810 102.310 138.855 ;
        RECT 104.800 138.810 105.090 138.855 ;
        RECT 106.660 138.810 106.950 138.855 ;
        RECT 102.020 138.670 106.950 138.810 ;
        RECT 102.020 138.625 102.310 138.670 ;
        RECT 104.800 138.625 105.090 138.670 ;
        RECT 106.660 138.625 106.950 138.670 ;
        RECT 61.200 138.330 68.240 138.470 ;
        RECT 47.770 138.270 48.090 138.330 ;
        RECT 50.070 138.270 50.390 138.330 ;
        RECT 53.750 138.270 54.070 138.330 ;
        RECT 66.630 138.270 66.950 138.330 ;
        RECT 79.510 138.270 79.830 138.530 ;
        RECT 90.105 138.470 90.395 138.515 ;
        RECT 91.010 138.470 91.330 138.530 ;
        RECT 90.105 138.330 91.330 138.470 ;
        RECT 90.105 138.285 90.395 138.330 ;
        RECT 91.010 138.270 91.330 138.330 ;
        RECT 98.370 138.470 98.690 138.530 ;
        RECT 107.200 138.470 107.340 138.965 ;
        RECT 110.420 138.810 110.560 139.340 ;
        RECT 110.805 139.320 111.095 139.340 ;
        RECT 111.265 139.305 111.555 139.535 ;
        RECT 111.725 139.305 112.015 139.535 ;
        RECT 111.340 139.150 111.480 139.305 ;
        RECT 112.630 139.290 112.950 139.550 ;
        RECT 112.720 139.150 112.860 139.290 ;
        RECT 111.340 139.010 112.860 139.150 ;
        RECT 112.630 138.810 112.950 138.870 ;
        RECT 114.100 138.810 114.240 139.690 ;
        RECT 117.015 139.645 117.550 139.690 ;
        RECT 119.020 139.830 119.310 139.875 ;
        RECT 120.450 139.830 120.770 139.890 ;
        RECT 122.280 139.830 122.570 139.875 ;
        RECT 119.020 139.690 122.570 139.830 ;
        RECT 119.020 139.645 119.310 139.690 ;
        RECT 117.230 139.630 117.550 139.645 ;
        RECT 120.450 139.630 120.770 139.690 ;
        RECT 122.280 139.645 122.570 139.690 ;
        RECT 123.200 139.830 123.490 139.875 ;
        RECT 125.060 139.830 125.350 139.875 ;
        RECT 123.200 139.690 125.350 139.830 ;
        RECT 123.200 139.645 123.490 139.690 ;
        RECT 125.060 139.645 125.350 139.690 ;
        RECT 115.405 139.305 115.695 139.535 ;
        RECT 110.420 138.670 114.240 138.810 ;
        RECT 115.480 138.810 115.620 139.305 ;
        RECT 115.850 139.290 116.170 139.550 ;
        RECT 120.880 139.490 121.170 139.535 ;
        RECT 123.200 139.490 123.415 139.645 ;
        RECT 120.880 139.350 123.415 139.490 ;
        RECT 120.880 139.305 121.170 139.350 ;
        RECT 124.130 139.290 124.450 139.550 ;
        RECT 125.970 138.950 126.290 139.210 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 119.990 138.810 120.310 138.870 ;
        RECT 115.480 138.670 120.310 138.810 ;
        RECT 112.630 138.610 112.950 138.670 ;
        RECT 119.990 138.610 120.310 138.670 ;
        RECT 120.880 138.810 121.170 138.855 ;
        RECT 123.660 138.810 123.950 138.855 ;
        RECT 125.520 138.810 125.810 138.855 ;
        RECT 120.880 138.670 125.810 138.810 ;
        RECT 120.880 138.625 121.170 138.670 ;
        RECT 123.660 138.625 123.950 138.670 ;
        RECT 125.520 138.625 125.810 138.670 ;
        RECT 121.370 138.470 121.690 138.530 ;
        RECT 124.590 138.470 124.910 138.530 ;
        RECT 126.060 138.470 126.200 138.950 ;
        RECT 98.370 138.330 126.200 138.470 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 98.370 138.270 98.690 138.330 ;
        RECT 121.370 138.270 121.690 138.330 ;
        RECT 124.590 138.270 124.910 138.330 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 14.580 137.650 127.740 138.130 ;
        RECT 34.430 137.250 34.750 137.510 ;
        RECT 35.825 137.265 36.115 137.495 ;
        RECT 38.110 137.450 38.430 137.510 ;
        RECT 38.585 137.450 38.875 137.495 ;
        RECT 38.110 137.310 38.875 137.450 ;
        RECT 33.970 137.110 34.290 137.170 ;
        RECT 35.900 137.110 36.040 137.265 ;
        RECT 38.110 137.250 38.430 137.310 ;
        RECT 38.585 137.265 38.875 137.310 ;
        RECT 44.550 137.250 44.870 137.510 ;
        RECT 48.230 137.450 48.550 137.510 ;
        RECT 50.990 137.450 51.310 137.510 ;
        RECT 53.290 137.450 53.610 137.510 ;
        RECT 48.230 137.310 53.610 137.450 ;
        RECT 48.230 137.250 48.550 137.310 ;
        RECT 50.990 137.250 51.310 137.310 ;
        RECT 53.290 137.250 53.610 137.310 ;
        RECT 60.650 137.450 60.970 137.510 ;
        RECT 60.650 137.310 62.720 137.450 ;
        RECT 60.650 137.250 60.970 137.310 ;
        RECT 61.125 137.110 61.415 137.155 ;
        RECT 33.970 136.970 36.040 137.110 ;
        RECT 40.040 136.970 61.415 137.110 ;
        RECT 33.970 136.910 34.290 136.970 ;
        RECT 21.550 136.770 21.870 136.830 ;
        RECT 22.945 136.770 23.235 136.815 ;
        RECT 21.550 136.630 23.235 136.770 ;
        RECT 21.550 136.570 21.870 136.630 ;
        RECT 22.945 136.585 23.235 136.630 ;
        RECT 31.210 136.570 31.530 136.830 ;
        RECT 35.350 136.770 35.670 136.830 ;
        RECT 36.285 136.770 36.575 136.815 ;
        RECT 35.350 136.630 36.575 136.770 ;
        RECT 35.350 136.570 35.670 136.630 ;
        RECT 36.285 136.585 36.575 136.630 ;
        RECT 39.030 136.570 39.350 136.830 ;
        RECT 22.025 136.430 22.315 136.475 ;
        RECT 22.470 136.430 22.790 136.490 ;
        RECT 22.025 136.290 22.790 136.430 ;
        RECT 22.025 136.245 22.315 136.290 ;
        RECT 22.470 136.230 22.790 136.290 ;
        RECT 32.605 136.245 32.895 136.475 ;
        RECT 33.510 136.430 33.830 136.490 ;
        RECT 34.890 136.430 35.210 136.490 ;
        RECT 33.510 136.290 35.210 136.430 ;
        RECT 30.290 136.090 30.610 136.150 ;
        RECT 22.560 135.950 30.610 136.090 ;
        RECT 18.790 135.750 19.110 135.810 ;
        RECT 20.185 135.750 20.475 135.795 ;
        RECT 18.790 135.610 20.475 135.750 ;
        RECT 18.790 135.550 19.110 135.610 ;
        RECT 20.185 135.565 20.475 135.610 ;
        RECT 22.010 135.750 22.330 135.810 ;
        RECT 22.560 135.795 22.700 135.950 ;
        RECT 30.290 135.890 30.610 135.950 ;
        RECT 32.680 135.810 32.820 136.245 ;
        RECT 33.510 136.230 33.830 136.290 ;
        RECT 34.890 136.230 35.210 136.290 ;
        RECT 35.825 136.430 36.115 136.475 ;
        RECT 36.730 136.430 37.050 136.490 ;
        RECT 35.825 136.290 37.050 136.430 ;
        RECT 35.825 136.245 36.115 136.290 ;
        RECT 36.730 136.230 37.050 136.290 ;
        RECT 38.570 136.230 38.890 136.490 ;
        RECT 40.040 136.475 40.180 136.970 ;
        RECT 61.125 136.925 61.415 136.970 ;
        RECT 62.580 137.110 62.720 137.310 ;
        RECT 65.250 137.250 65.570 137.510 ;
        RECT 71.245 137.450 71.535 137.495 ;
        RECT 74.910 137.450 75.230 137.510 ;
        RECT 71.245 137.310 75.230 137.450 ;
        RECT 71.245 137.265 71.535 137.310 ;
        RECT 74.910 137.250 75.230 137.310 ;
        RECT 79.525 137.450 79.815 137.495 ;
        RECT 79.970 137.450 80.290 137.510 ;
        RECT 83.895 137.450 84.185 137.495 ;
        RECT 84.570 137.450 84.890 137.510 ;
        RECT 79.525 137.310 80.290 137.450 ;
        RECT 79.525 137.265 79.815 137.310 ;
        RECT 79.970 137.250 80.290 137.310 ;
        RECT 81.440 137.310 82.960 137.450 ;
        RECT 65.340 137.110 65.480 137.250 ;
        RECT 74.450 137.110 74.770 137.170 ;
        RECT 62.580 136.970 74.770 137.110 ;
        RECT 45.470 136.570 45.790 136.830 ;
        RECT 50.530 136.770 50.850 136.830 ;
        RECT 48.780 136.630 50.850 136.770 ;
        RECT 39.965 136.245 40.255 136.475 ;
        RECT 42.250 136.430 42.570 136.490 ;
        RECT 44.565 136.430 44.855 136.475 ;
        RECT 42.250 136.290 44.855 136.430 ;
        RECT 42.250 136.230 42.570 136.290 ;
        RECT 44.565 136.245 44.855 136.290 ;
        RECT 45.560 136.290 47.540 136.430 ;
        RECT 37.205 136.090 37.495 136.135 ;
        RECT 45.560 136.090 45.700 136.290 ;
        RECT 37.205 135.950 45.700 136.090 ;
        RECT 45.945 136.090 46.235 136.135 ;
        RECT 46.405 136.090 46.695 136.135 ;
        RECT 45.945 135.950 46.695 136.090 ;
        RECT 47.400 136.090 47.540 136.290 ;
        RECT 47.770 136.230 48.090 136.490 ;
        RECT 48.230 136.230 48.550 136.490 ;
        RECT 48.780 136.475 48.920 136.630 ;
        RECT 50.530 136.570 50.850 136.630 ;
        RECT 54.225 136.770 54.515 136.815 ;
        RECT 54.670 136.770 54.990 136.830 ;
        RECT 54.225 136.630 54.990 136.770 ;
        RECT 54.225 136.585 54.515 136.630 ;
        RECT 54.670 136.570 54.990 136.630 ;
        RECT 48.705 136.245 48.995 136.475 ;
        RECT 49.625 136.245 49.915 136.475 ;
        RECT 50.620 136.430 50.760 136.570 ;
        RECT 62.580 136.475 62.720 136.970 ;
        RECT 74.450 136.910 74.770 136.970 ;
        RECT 77.225 137.110 77.515 137.155 ;
        RECT 81.440 137.110 81.580 137.310 ;
        RECT 82.270 137.110 82.590 137.170 ;
        RECT 77.225 136.970 81.580 137.110 ;
        RECT 81.900 136.970 82.590 137.110 ;
        RECT 82.820 137.110 82.960 137.310 ;
        RECT 83.895 137.310 84.890 137.450 ;
        RECT 83.895 137.265 84.185 137.310 ;
        RECT 84.570 137.250 84.890 137.310 ;
        RECT 85.030 137.450 85.350 137.510 ;
        RECT 105.270 137.450 105.590 137.510 ;
        RECT 107.125 137.450 107.415 137.495 ;
        RECT 85.030 137.310 95.840 137.450 ;
        RECT 85.030 137.250 85.350 137.310 ;
        RECT 86.870 137.110 87.190 137.170 ;
        RECT 82.820 136.970 87.190 137.110 ;
        RECT 77.225 136.925 77.515 136.970 ;
        RECT 65.265 136.770 65.555 136.815 ;
        RECT 65.710 136.770 66.030 136.830 ;
        RECT 73.990 136.770 74.310 136.830 ;
        RECT 63.040 136.630 64.100 136.770 ;
        RECT 63.040 136.475 63.180 136.630 ;
        RECT 55.145 136.430 55.435 136.475 ;
        RECT 57.905 136.430 58.195 136.475 ;
        RECT 50.620 136.290 55.435 136.430 ;
        RECT 55.145 136.245 55.435 136.290 ;
        RECT 57.060 136.290 58.195 136.430 ;
        RECT 49.150 136.090 49.470 136.150 ;
        RECT 47.400 135.950 49.470 136.090 ;
        RECT 49.700 136.090 49.840 136.245 ;
        RECT 50.530 136.090 50.850 136.150 ;
        RECT 52.370 136.090 52.690 136.150 ;
        RECT 55.590 136.090 55.910 136.150 ;
        RECT 49.700 135.950 55.910 136.090 ;
        RECT 37.205 135.905 37.495 135.950 ;
        RECT 45.945 135.905 46.235 135.950 ;
        RECT 46.405 135.905 46.695 135.950 ;
        RECT 49.150 135.890 49.470 135.950 ;
        RECT 50.530 135.890 50.850 135.950 ;
        RECT 52.370 135.890 52.690 135.950 ;
        RECT 55.590 135.890 55.910 135.950 ;
        RECT 22.485 135.750 22.775 135.795 ;
        RECT 22.010 135.610 22.775 135.750 ;
        RECT 22.010 135.550 22.330 135.610 ;
        RECT 22.485 135.565 22.775 135.610 ;
        RECT 28.450 135.550 28.770 135.810 ;
        RECT 30.750 135.750 31.070 135.810 ;
        RECT 32.590 135.750 32.910 135.810 ;
        RECT 30.750 135.610 32.910 135.750 ;
        RECT 30.750 135.550 31.070 135.610 ;
        RECT 32.590 135.550 32.910 135.610 ;
        RECT 34.430 135.750 34.750 135.810 ;
        RECT 34.905 135.750 35.195 135.795 ;
        RECT 34.430 135.610 35.195 135.750 ;
        RECT 34.430 135.550 34.750 135.610 ;
        RECT 34.905 135.565 35.195 135.610 ;
        RECT 37.665 135.750 37.955 135.795 ;
        RECT 38.570 135.750 38.890 135.810 ;
        RECT 37.665 135.610 38.890 135.750 ;
        RECT 37.665 135.565 37.955 135.610 ;
        RECT 38.570 135.550 38.890 135.610 ;
        RECT 43.645 135.750 43.935 135.795 ;
        RECT 51.910 135.750 52.230 135.810 ;
        RECT 43.645 135.610 52.230 135.750 ;
        RECT 43.645 135.565 43.935 135.610 ;
        RECT 51.910 135.550 52.230 135.610 ;
        RECT 54.685 135.750 54.975 135.795 ;
        RECT 56.510 135.750 56.830 135.810 ;
        RECT 57.060 135.795 57.200 136.290 ;
        RECT 57.905 136.245 58.195 136.290 ;
        RECT 62.505 136.245 62.795 136.475 ;
        RECT 62.965 136.245 63.255 136.475 ;
        RECT 63.425 136.245 63.715 136.475 ;
        RECT 60.650 136.090 60.970 136.150 ;
        RECT 63.500 136.090 63.640 136.245 ;
        RECT 60.650 135.950 63.640 136.090 ;
        RECT 63.960 136.090 64.100 136.630 ;
        RECT 65.265 136.630 66.030 136.770 ;
        RECT 65.265 136.585 65.555 136.630 ;
        RECT 65.710 136.570 66.030 136.630 ;
        RECT 69.940 136.630 74.310 136.770 ;
        RECT 64.330 136.230 64.650 136.490 ;
        RECT 68.025 136.430 68.315 136.475 ;
        RECT 68.485 136.430 68.775 136.475 ;
        RECT 68.025 136.290 68.775 136.430 ;
        RECT 68.025 136.245 68.315 136.290 ;
        RECT 68.485 136.245 68.775 136.290 ;
        RECT 69.390 136.230 69.710 136.490 ;
        RECT 69.940 136.475 70.080 136.630 ;
        RECT 73.990 136.570 74.310 136.630 ;
        RECT 69.865 136.245 70.155 136.475 ;
        RECT 70.325 136.245 70.615 136.475 ;
        RECT 76.290 136.430 76.610 136.490 ;
        RECT 78.145 136.430 78.435 136.475 ;
        RECT 76.290 136.290 78.435 136.430 ;
        RECT 65.250 136.090 65.570 136.150 ;
        RECT 66.630 136.090 66.950 136.150 ;
        RECT 70.400 136.090 70.540 136.245 ;
        RECT 76.290 136.230 76.610 136.290 ;
        RECT 78.145 136.245 78.435 136.290 ;
        RECT 78.605 136.245 78.895 136.475 ;
        RECT 63.960 135.950 66.950 136.090 ;
        RECT 60.650 135.890 60.970 135.950 ;
        RECT 65.250 135.890 65.570 135.950 ;
        RECT 66.630 135.890 66.950 135.950 ;
        RECT 69.940 135.950 70.540 136.090 ;
        RECT 78.680 136.090 78.820 136.245 ;
        RECT 79.510 136.230 79.830 136.490 ;
        RECT 81.350 136.230 81.670 136.490 ;
        RECT 81.900 136.475 82.040 136.970 ;
        RECT 82.270 136.910 82.590 136.970 ;
        RECT 86.870 136.910 87.190 136.970 ;
        RECT 87.760 137.110 88.050 137.155 ;
        RECT 90.540 137.110 90.830 137.155 ;
        RECT 92.400 137.110 92.690 137.155 ;
        RECT 87.760 136.970 92.690 137.110 ;
        RECT 95.700 137.110 95.840 137.310 ;
        RECT 105.270 137.310 107.415 137.450 ;
        RECT 105.270 137.250 105.590 137.310 ;
        RECT 107.125 137.265 107.415 137.310 ;
        RECT 119.530 137.450 119.850 137.510 ;
        RECT 119.530 137.310 123.440 137.450 ;
        RECT 119.530 137.250 119.850 137.310 ;
        RECT 113.090 137.110 113.410 137.170 ;
        RECT 95.700 136.970 96.300 137.110 ;
        RECT 87.760 136.925 88.050 136.970 ;
        RECT 90.540 136.925 90.830 136.970 ;
        RECT 92.400 136.925 92.690 136.970 ;
        RECT 86.410 136.770 86.730 136.830 ;
        RECT 82.360 136.630 86.730 136.770 ;
        RECT 82.360 136.475 82.500 136.630 ;
        RECT 86.410 136.570 86.730 136.630 ;
        RECT 91.010 136.570 91.330 136.830 ;
        RECT 91.470 136.770 91.790 136.830 ;
        RECT 96.160 136.815 96.300 136.970 ;
        RECT 103.520 136.970 113.410 137.110 ;
        RECT 103.520 136.815 103.660 136.970 ;
        RECT 109.960 136.815 110.100 136.970 ;
        RECT 113.090 136.910 113.410 136.970 ;
        RECT 117.660 137.110 117.950 137.155 ;
        RECT 120.440 137.110 120.730 137.155 ;
        RECT 122.300 137.110 122.590 137.155 ;
        RECT 117.660 136.970 122.590 137.110 ;
        RECT 117.660 136.925 117.950 136.970 ;
        RECT 120.440 136.925 120.730 136.970 ;
        RECT 122.300 136.925 122.590 136.970 ;
        RECT 95.625 136.770 95.915 136.815 ;
        RECT 91.470 136.630 95.915 136.770 ;
        RECT 91.470 136.570 91.790 136.630 ;
        RECT 95.625 136.585 95.915 136.630 ;
        RECT 96.085 136.770 96.375 136.815 ;
        RECT 103.445 136.770 103.735 136.815 ;
        RECT 96.085 136.630 103.735 136.770 ;
        RECT 96.085 136.585 96.375 136.630 ;
        RECT 103.445 136.585 103.735 136.630 ;
        RECT 104.900 136.630 109.180 136.770 ;
        RECT 81.825 136.245 82.115 136.475 ;
        RECT 82.285 136.245 82.575 136.475 ;
        RECT 83.190 136.230 83.510 136.490 ;
        RECT 87.760 136.430 88.050 136.475 ;
        RECT 87.760 136.290 90.295 136.430 ;
        RECT 87.760 136.245 88.050 136.290 ;
        RECT 84.110 136.090 84.430 136.150 ;
        RECT 78.680 135.950 84.430 136.090 ;
        RECT 54.685 135.610 56.830 135.750 ;
        RECT 54.685 135.565 54.975 135.610 ;
        RECT 56.510 135.550 56.830 135.610 ;
        RECT 56.985 135.565 57.275 135.795 ;
        RECT 58.825 135.750 59.115 135.795 ;
        RECT 59.730 135.750 60.050 135.810 ;
        RECT 58.825 135.610 60.050 135.750 ;
        RECT 58.825 135.565 59.115 135.610 ;
        RECT 59.730 135.550 60.050 135.610 ;
        RECT 61.110 135.750 61.430 135.810 ;
        RECT 69.940 135.750 70.080 135.950 ;
        RECT 84.110 135.890 84.430 135.950 ;
        RECT 85.900 136.090 86.190 136.135 ;
        RECT 88.250 136.090 88.570 136.150 ;
        RECT 90.080 136.135 90.295 136.290 ;
        RECT 92.865 136.245 93.155 136.475 ;
        RECT 93.310 136.430 93.630 136.490 ;
        RECT 97.910 136.430 98.230 136.490 ;
        RECT 93.310 136.290 98.230 136.430 ;
        RECT 89.160 136.090 89.450 136.135 ;
        RECT 85.900 135.950 89.450 136.090 ;
        RECT 85.900 135.905 86.190 135.950 ;
        RECT 88.250 135.890 88.570 135.950 ;
        RECT 89.160 135.905 89.450 135.950 ;
        RECT 90.080 136.090 90.370 136.135 ;
        RECT 91.940 136.090 92.230 136.135 ;
        RECT 90.080 135.950 92.230 136.090 ;
        RECT 92.940 136.090 93.080 136.245 ;
        RECT 93.310 136.230 93.630 136.290 ;
        RECT 97.910 136.230 98.230 136.290 ;
        RECT 98.830 136.230 99.150 136.490 ;
        RECT 99.290 136.230 99.610 136.490 ;
        RECT 99.765 136.430 100.055 136.475 ;
        RECT 100.210 136.430 100.530 136.490 ;
        RECT 104.900 136.475 105.040 136.630 ;
        RECT 104.365 136.430 104.655 136.475 ;
        RECT 99.765 136.290 100.530 136.430 ;
        RECT 99.765 136.245 100.055 136.290 ;
        RECT 100.210 136.230 100.530 136.290 ;
        RECT 100.760 136.290 104.655 136.430 ;
        RECT 94.230 136.090 94.550 136.150 ;
        RECT 98.370 136.090 98.690 136.150 ;
        RECT 92.940 135.950 98.690 136.090 ;
        RECT 90.080 135.905 90.370 135.950 ;
        RECT 91.940 135.905 92.230 135.950 ;
        RECT 94.230 135.890 94.550 135.950 ;
        RECT 98.370 135.890 98.690 135.950 ;
        RECT 98.920 136.090 99.060 136.230 ;
        RECT 100.760 136.090 100.900 136.290 ;
        RECT 104.365 136.245 104.655 136.290 ;
        RECT 104.825 136.245 105.115 136.475 ;
        RECT 108.045 136.430 108.335 136.475 ;
        RECT 106.740 136.290 108.335 136.430 ;
        RECT 98.920 135.950 100.900 136.090 ;
        RECT 61.110 135.610 70.080 135.750 ;
        RECT 79.050 135.750 79.370 135.810 ;
        RECT 79.985 135.750 80.275 135.795 ;
        RECT 79.050 135.610 80.275 135.750 ;
        RECT 61.110 135.550 61.430 135.610 ;
        RECT 79.050 135.550 79.370 135.610 ;
        RECT 79.985 135.565 80.275 135.610 ;
        RECT 85.030 135.750 85.350 135.810 ;
        RECT 92.850 135.750 93.170 135.810 ;
        RECT 85.030 135.610 93.170 135.750 ;
        RECT 85.030 135.550 85.350 135.610 ;
        RECT 92.850 135.550 93.170 135.610 ;
        RECT 93.325 135.750 93.615 135.795 ;
        RECT 93.770 135.750 94.090 135.810 ;
        RECT 93.325 135.610 94.090 135.750 ;
        RECT 93.325 135.565 93.615 135.610 ;
        RECT 93.770 135.550 94.090 135.610 ;
        RECT 95.165 135.750 95.455 135.795 ;
        RECT 98.920 135.750 99.060 135.950 ;
        RECT 95.165 135.610 99.060 135.750 ;
        RECT 95.165 135.565 95.455 135.610 ;
        RECT 101.130 135.550 101.450 135.810 ;
        RECT 106.740 135.795 106.880 136.290 ;
        RECT 108.045 136.245 108.335 136.290 ;
        RECT 109.040 136.150 109.180 136.630 ;
        RECT 109.885 136.585 110.175 136.815 ;
        RECT 121.370 136.770 121.690 136.830 ;
        RECT 122.765 136.770 123.055 136.815 ;
        RECT 121.370 136.630 123.055 136.770 ;
        RECT 121.370 136.570 121.690 136.630 ;
        RECT 122.765 136.585 123.055 136.630 ;
        RECT 111.265 136.430 111.555 136.475 ;
        RECT 112.630 136.430 112.950 136.490 ;
        RECT 111.265 136.290 112.950 136.430 ;
        RECT 111.265 136.245 111.555 136.290 ;
        RECT 112.630 136.230 112.950 136.290 ;
        RECT 117.660 136.430 117.950 136.475 ;
        RECT 117.660 136.290 120.195 136.430 ;
        RECT 117.660 136.245 117.950 136.290 ;
        RECT 108.950 136.090 109.270 136.150 ;
        RECT 115.850 136.135 116.170 136.150 ;
        RECT 119.980 136.135 120.195 136.290 ;
        RECT 120.910 136.230 121.230 136.490 ;
        RECT 123.300 136.475 123.440 137.310 ;
        RECT 124.130 137.250 124.450 137.510 ;
        RECT 123.225 136.245 123.515 136.475 ;
        RECT 110.805 136.090 111.095 136.135 ;
        RECT 113.795 136.090 114.085 136.135 ;
        RECT 108.950 135.950 114.085 136.090 ;
        RECT 108.950 135.890 109.270 135.950 ;
        RECT 110.805 135.905 111.095 135.950 ;
        RECT 113.795 135.905 114.085 135.950 ;
        RECT 115.800 136.090 116.170 136.135 ;
        RECT 119.060 136.090 119.350 136.135 ;
        RECT 115.800 135.950 119.350 136.090 ;
        RECT 115.800 135.905 116.170 135.950 ;
        RECT 119.060 135.905 119.350 135.950 ;
        RECT 119.980 136.090 120.270 136.135 ;
        RECT 121.840 136.090 122.130 136.135 ;
        RECT 119.980 135.950 122.130 136.090 ;
        RECT 119.980 135.905 120.270 135.950 ;
        RECT 121.840 135.905 122.130 135.950 ;
        RECT 115.850 135.890 116.170 135.905 ;
        RECT 106.665 135.565 106.955 135.795 ;
        RECT 113.090 135.550 113.410 135.810 ;
        RECT 14.580 134.930 127.740 135.410 ;
        RECT 19.250 134.530 19.570 134.790 ;
        RECT 20.875 134.730 21.165 134.775 ;
        RECT 22.010 134.730 22.330 134.790 ;
        RECT 20.875 134.590 22.330 134.730 ;
        RECT 20.875 134.545 21.165 134.590 ;
        RECT 22.010 134.530 22.330 134.590 ;
        RECT 32.605 134.730 32.895 134.775 ;
        RECT 33.970 134.730 34.290 134.790 ;
        RECT 32.605 134.590 34.290 134.730 ;
        RECT 32.605 134.545 32.895 134.590 ;
        RECT 33.970 134.530 34.290 134.590 ;
        RECT 50.530 134.530 50.850 134.790 ;
        RECT 52.615 134.730 52.905 134.775 ;
        RECT 56.510 134.730 56.830 134.790 ;
        RECT 51.080 134.590 56.830 134.730 ;
        RECT 16.965 134.390 17.255 134.435 ;
        RECT 19.340 134.390 19.480 134.530 ;
        RECT 16.965 134.250 19.480 134.390 ;
        RECT 19.725 134.390 20.015 134.435 ;
        RECT 22.880 134.390 23.170 134.435 ;
        RECT 26.140 134.390 26.430 134.435 ;
        RECT 19.725 134.250 26.430 134.390 ;
        RECT 16.965 134.205 17.255 134.250 ;
        RECT 19.725 134.205 20.015 134.250 ;
        RECT 22.880 134.205 23.170 134.250 ;
        RECT 26.140 134.205 26.430 134.250 ;
        RECT 27.060 134.390 27.350 134.435 ;
        RECT 28.920 134.390 29.210 134.435 ;
        RECT 36.270 134.390 36.590 134.450 ;
        RECT 27.060 134.250 29.210 134.390 ;
        RECT 27.060 134.205 27.350 134.250 ;
        RECT 28.920 134.205 29.210 134.250 ;
        RECT 29.920 134.250 36.590 134.390 ;
        RECT 17.425 133.865 17.715 134.095 ;
        RECT 17.885 134.050 18.175 134.095 ;
        RECT 18.790 134.050 19.110 134.110 ;
        RECT 17.885 133.910 19.110 134.050 ;
        RECT 17.885 133.865 18.175 133.910 ;
        RECT 17.500 133.710 17.640 133.865 ;
        RECT 18.790 133.850 19.110 133.910 ;
        RECT 19.265 134.050 19.555 134.095 ;
        RECT 24.740 134.050 25.030 134.095 ;
        RECT 27.060 134.050 27.275 134.205 ;
        RECT 29.920 134.110 30.060 134.250 ;
        RECT 36.270 134.190 36.590 134.250 ;
        RECT 42.265 134.390 42.555 134.435 ;
        RECT 48.705 134.390 48.995 134.435 ;
        RECT 50.620 134.390 50.760 134.530 ;
        RECT 42.265 134.250 48.995 134.390 ;
        RECT 42.265 134.205 42.555 134.250 ;
        RECT 48.705 134.205 48.995 134.250 ;
        RECT 49.700 134.250 50.760 134.390 ;
        RECT 19.265 133.910 19.940 134.050 ;
        RECT 19.265 133.865 19.555 133.910 ;
        RECT 19.800 133.770 19.940 133.910 ;
        RECT 24.740 133.910 27.275 134.050 ;
        RECT 27.620 133.910 29.600 134.050 ;
        RECT 24.740 133.865 25.030 133.910 ;
        RECT 19.710 133.710 20.030 133.770 ;
        RECT 17.500 133.570 20.030 133.710 ;
        RECT 19.710 133.510 20.030 133.570 ;
        RECT 22.010 133.710 22.330 133.770 ;
        RECT 27.620 133.710 27.760 133.910 ;
        RECT 22.010 133.570 27.760 133.710 ;
        RECT 28.005 133.710 28.295 133.755 ;
        RECT 28.910 133.710 29.230 133.770 ;
        RECT 28.005 133.570 29.230 133.710 ;
        RECT 29.460 133.710 29.600 133.910 ;
        RECT 29.830 133.850 30.150 134.110 ;
        RECT 31.210 134.050 31.530 134.110 ;
        RECT 30.380 133.910 31.530 134.050 ;
        RECT 30.380 133.710 30.520 133.910 ;
        RECT 31.210 133.850 31.530 133.910 ;
        RECT 31.685 134.050 31.975 134.095 ;
        RECT 32.130 134.050 32.450 134.110 ;
        RECT 31.685 133.910 32.450 134.050 ;
        RECT 31.685 133.865 31.975 133.910 ;
        RECT 32.130 133.850 32.450 133.910 ;
        RECT 32.590 134.050 32.910 134.110 ;
        RECT 34.905 134.050 35.195 134.095 ;
        RECT 32.590 133.910 35.195 134.050 ;
        RECT 32.590 133.850 32.910 133.910 ;
        RECT 34.905 133.865 35.195 133.910 ;
        RECT 39.505 133.865 39.795 134.095 ;
        RECT 29.460 133.570 30.520 133.710 ;
        RECT 22.010 133.510 22.330 133.570 ;
        RECT 28.005 133.525 28.295 133.570 ;
        RECT 28.910 133.510 29.230 133.570 ;
        RECT 30.765 133.525 31.055 133.755 ;
        RECT 31.300 133.710 31.440 133.850 ;
        RECT 33.525 133.710 33.815 133.755 ;
        RECT 31.300 133.570 33.815 133.710 ;
        RECT 33.525 133.525 33.815 133.570 ;
        RECT 34.445 133.525 34.735 133.755 ;
        RECT 39.580 133.710 39.720 133.865 ;
        RECT 40.410 133.850 40.730 134.110 ;
        RECT 40.870 133.850 41.190 134.110 ;
        RECT 42.710 134.050 43.030 134.110 ;
        RECT 43.185 134.050 43.475 134.095 ;
        RECT 42.710 133.910 43.475 134.050 ;
        RECT 42.710 133.850 43.030 133.910 ;
        RECT 43.185 133.865 43.475 133.910 ;
        RECT 43.630 133.850 43.950 134.110 ;
        RECT 46.390 133.850 46.710 134.110 ;
        RECT 46.865 133.865 47.155 134.095 ;
        RECT 47.325 133.865 47.615 134.095 ;
        RECT 48.245 134.050 48.535 134.095 ;
        RECT 49.700 134.050 49.840 134.250 ;
        RECT 48.245 133.910 49.840 134.050 ;
        RECT 48.245 133.865 48.535 133.910 ;
        RECT 45.025 133.710 45.315 133.755 ;
        RECT 39.580 133.570 45.315 133.710 ;
        RECT 45.025 133.525 45.315 133.570 ;
        RECT 18.805 133.370 19.095 133.415 ;
        RECT 23.390 133.370 23.710 133.430 ;
        RECT 18.805 133.230 23.710 133.370 ;
        RECT 18.805 133.185 19.095 133.230 ;
        RECT 23.390 133.170 23.710 133.230 ;
        RECT 24.740 133.370 25.030 133.415 ;
        RECT 27.520 133.370 27.810 133.415 ;
        RECT 29.380 133.370 29.670 133.415 ;
        RECT 24.740 133.230 29.670 133.370 ;
        RECT 30.840 133.370 30.980 133.525 ;
        RECT 34.520 133.370 34.660 133.525 ;
        RECT 34.890 133.370 35.210 133.430 ;
        RECT 30.840 133.230 35.210 133.370 ;
        RECT 24.740 133.185 25.030 133.230 ;
        RECT 27.520 133.185 27.810 133.230 ;
        RECT 29.380 133.185 29.670 133.230 ;
        RECT 34.890 133.170 35.210 133.230 ;
        RECT 31.210 133.030 31.530 133.090 ;
        RECT 35.810 133.030 36.130 133.090 ;
        RECT 31.210 132.890 36.130 133.030 ;
        RECT 31.210 132.830 31.530 132.890 ;
        RECT 35.810 132.830 36.130 132.890 ;
        RECT 36.745 133.030 37.035 133.075 ;
        RECT 39.490 133.030 39.810 133.090 ;
        RECT 36.745 132.890 39.810 133.030 ;
        RECT 36.745 132.845 37.035 132.890 ;
        RECT 39.490 132.830 39.810 132.890 ;
        RECT 40.410 132.830 40.730 133.090 ;
        RECT 41.330 133.030 41.650 133.090 ;
        RECT 41.805 133.030 42.095 133.075 ;
        RECT 41.330 132.890 42.095 133.030 ;
        RECT 41.330 132.830 41.650 132.890 ;
        RECT 41.805 132.845 42.095 132.890 ;
        RECT 43.170 132.830 43.490 133.090 ;
        RECT 44.090 133.030 44.410 133.090 ;
        RECT 44.565 133.030 44.855 133.075 ;
        RECT 44.090 132.890 44.855 133.030 ;
        RECT 46.940 133.030 47.080 133.865 ;
        RECT 47.400 133.370 47.540 133.865 ;
        RECT 50.070 133.850 50.390 134.110 ;
        RECT 50.530 133.850 50.850 134.110 ;
        RECT 51.080 134.095 51.220 134.590 ;
        RECT 52.615 134.545 52.905 134.590 ;
        RECT 56.510 134.530 56.830 134.590 ;
        RECT 74.450 134.730 74.770 134.790 ;
        RECT 87.805 134.730 88.095 134.775 ;
        RECT 88.250 134.730 88.570 134.790 ;
        RECT 100.210 134.730 100.530 134.790 ;
        RECT 102.065 134.730 102.355 134.775 ;
        RECT 102.510 134.730 102.830 134.790 ;
        RECT 74.450 134.590 87.560 134.730 ;
        RECT 74.450 134.530 74.770 134.590 ;
        RECT 54.620 134.390 54.910 134.435 ;
        RECT 56.050 134.390 56.370 134.450 ;
        RECT 57.880 134.390 58.170 134.435 ;
        RECT 54.620 134.250 58.170 134.390 ;
        RECT 54.620 134.205 54.910 134.250 ;
        RECT 56.050 134.190 56.370 134.250 ;
        RECT 57.880 134.205 58.170 134.250 ;
        RECT 58.800 134.390 59.090 134.435 ;
        RECT 60.660 134.390 60.950 134.435 ;
        RECT 58.800 134.250 60.950 134.390 ;
        RECT 58.800 134.205 59.090 134.250 ;
        RECT 60.660 134.205 60.950 134.250 ;
        RECT 64.330 134.390 64.650 134.450 ;
        RECT 64.330 134.250 66.860 134.390 ;
        RECT 51.005 133.865 51.295 134.095 ;
        RECT 51.925 134.050 52.215 134.095 ;
        RECT 52.370 134.050 52.690 134.110 ;
        RECT 51.925 133.910 52.690 134.050 ;
        RECT 51.925 133.865 52.215 133.910 ;
        RECT 52.370 133.850 52.690 133.910 ;
        RECT 56.480 134.050 56.770 134.095 ;
        RECT 58.800 134.050 59.015 134.205 ;
        RECT 64.330 134.190 64.650 134.250 ;
        RECT 56.480 133.910 59.015 134.050 ;
        RECT 56.480 133.865 56.770 133.910 ;
        RECT 59.730 133.850 60.050 134.110 ;
        RECT 61.585 134.050 61.875 134.095 ;
        RECT 63.870 134.050 64.190 134.110 ;
        RECT 61.585 133.910 64.190 134.050 ;
        RECT 61.585 133.865 61.875 133.910 ;
        RECT 63.870 133.850 64.190 133.910 ;
        RECT 64.790 133.850 65.110 134.110 ;
        RECT 65.250 133.850 65.570 134.110 ;
        RECT 65.710 133.850 66.030 134.110 ;
        RECT 66.720 134.095 66.860 134.250 ;
        RECT 79.050 134.190 79.370 134.450 ;
        RECT 85.030 134.390 85.350 134.450 ;
        RECT 80.060 134.250 85.350 134.390 ;
        RECT 87.420 134.390 87.560 134.590 ;
        RECT 87.805 134.590 88.570 134.730 ;
        RECT 87.805 134.545 88.095 134.590 ;
        RECT 88.250 134.530 88.570 134.590 ;
        RECT 90.180 134.590 101.820 134.730 ;
        RECT 90.180 134.390 90.320 134.590 ;
        RECT 100.210 134.530 100.530 134.590 ;
        RECT 87.420 134.250 90.320 134.390 ;
        RECT 90.550 134.390 90.870 134.450 ;
        RECT 91.420 134.390 91.710 134.435 ;
        RECT 94.680 134.390 94.970 134.435 ;
        RECT 90.550 134.250 94.970 134.390 ;
        RECT 66.645 134.050 66.935 134.095 ;
        RECT 80.060 134.050 80.200 134.250 ;
        RECT 85.030 134.190 85.350 134.250 ;
        RECT 90.550 134.190 90.870 134.250 ;
        RECT 91.420 134.205 91.710 134.250 ;
        RECT 94.680 134.205 94.970 134.250 ;
        RECT 95.600 134.390 95.890 134.435 ;
        RECT 97.460 134.390 97.750 134.435 ;
        RECT 95.600 134.250 97.750 134.390 ;
        RECT 95.600 134.205 95.890 134.250 ;
        RECT 97.460 134.205 97.750 134.250 ;
        RECT 66.645 133.910 80.200 134.050 ;
        RECT 66.645 133.865 66.935 133.910 ;
        RECT 80.430 133.850 80.750 134.110 ;
        RECT 88.250 133.850 88.570 134.110 ;
        RECT 93.280 134.050 93.570 134.095 ;
        RECT 95.600 134.050 95.815 134.205 ;
        RECT 101.130 134.190 101.450 134.450 ;
        RECT 101.680 134.390 101.820 134.590 ;
        RECT 102.065 134.590 102.830 134.730 ;
        RECT 102.065 134.545 102.355 134.590 ;
        RECT 102.510 134.530 102.830 134.590 ;
        RECT 120.005 134.730 120.295 134.775 ;
        RECT 120.910 134.730 121.230 134.790 ;
        RECT 120.005 134.590 121.230 134.730 ;
        RECT 120.005 134.545 120.295 134.590 ;
        RECT 120.910 134.530 121.230 134.590 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 105.745 134.390 106.035 134.435 ;
        RECT 106.205 134.390 106.495 134.435 ;
        RECT 110.330 134.390 110.650 134.450 ;
        RECT 101.680 134.250 104.940 134.390 ;
        RECT 93.280 133.910 95.815 134.050 ;
        RECT 93.280 133.865 93.570 133.910 ;
        RECT 97.910 133.850 98.230 134.110 ;
        RECT 98.370 133.850 98.690 134.110 ;
        RECT 99.750 133.850 100.070 134.110 ;
        RECT 102.510 133.850 102.830 134.110 ;
        RECT 103.890 134.050 104.210 134.110 ;
        RECT 104.365 134.050 104.655 134.095 ;
        RECT 103.890 133.910 104.655 134.050 ;
        RECT 104.800 134.050 104.940 134.250 ;
        RECT 105.745 134.250 106.495 134.390 ;
        RECT 105.745 134.205 106.035 134.250 ;
        RECT 106.205 134.205 106.495 134.250 ;
        RECT 107.660 134.250 110.650 134.390 ;
        RECT 107.660 134.095 107.800 134.250 ;
        RECT 110.330 134.190 110.650 134.250 ;
        RECT 112.170 134.190 112.490 134.450 ;
        RECT 107.585 134.050 107.875 134.095 ;
        RECT 104.800 133.910 107.875 134.050 ;
        RECT 103.890 133.850 104.210 133.910 ;
        RECT 104.365 133.865 104.655 133.910 ;
        RECT 107.585 133.865 107.875 133.910 ;
        RECT 108.030 133.850 108.350 134.110 ;
        RECT 108.505 134.050 108.795 134.095 ;
        RECT 108.950 134.050 109.270 134.110 ;
        RECT 108.505 133.910 109.270 134.050 ;
        RECT 108.505 133.865 108.795 133.910 ;
        RECT 108.950 133.850 109.270 133.910 ;
        RECT 109.410 133.850 109.730 134.110 ;
        RECT 110.790 133.850 111.110 134.110 ;
        RECT 111.250 133.850 111.570 134.110 ;
        RECT 113.090 134.050 113.410 134.110 ;
        RECT 119.085 134.050 119.375 134.095 ;
        RECT 113.090 133.910 119.375 134.050 ;
        RECT 113.090 133.850 113.410 133.910 ;
        RECT 119.085 133.865 119.375 133.910 ;
        RECT 49.150 133.710 49.470 133.770 ;
        RECT 63.425 133.710 63.715 133.755 ;
        RECT 49.150 133.570 63.715 133.710 ;
        RECT 49.150 133.510 49.470 133.570 ;
        RECT 63.425 133.525 63.715 133.570 ;
        RECT 79.985 133.710 80.275 133.755 ;
        RECT 83.650 133.710 83.970 133.770 ;
        RECT 79.985 133.570 83.970 133.710 ;
        RECT 79.985 133.525 80.275 133.570 ;
        RECT 83.650 133.510 83.970 133.570 ;
        RECT 86.410 133.710 86.730 133.770 ;
        RECT 89.415 133.710 89.705 133.755 ;
        RECT 91.470 133.710 91.790 133.770 ;
        RECT 86.410 133.570 91.790 133.710 ;
        RECT 86.410 133.510 86.730 133.570 ;
        RECT 89.415 133.525 89.705 133.570 ;
        RECT 91.470 133.510 91.790 133.570 ;
        RECT 95.150 133.710 95.470 133.770 ;
        RECT 96.545 133.710 96.835 133.755 ;
        RECT 95.150 133.570 96.835 133.710 ;
        RECT 98.000 133.710 98.140 133.850 ;
        RECT 98.000 133.570 100.440 133.710 ;
        RECT 95.150 133.510 95.470 133.570 ;
        RECT 96.545 133.525 96.835 133.570 ;
        RECT 55.590 133.370 55.910 133.430 ;
        RECT 47.400 133.230 55.910 133.370 ;
        RECT 55.590 133.170 55.910 133.230 ;
        RECT 56.480 133.370 56.770 133.415 ;
        RECT 59.260 133.370 59.550 133.415 ;
        RECT 61.120 133.370 61.410 133.415 ;
        RECT 56.480 133.230 61.410 133.370 ;
        RECT 56.480 133.185 56.770 133.230 ;
        RECT 59.260 133.185 59.550 133.230 ;
        RECT 61.120 133.185 61.410 133.230 ;
        RECT 81.365 133.370 81.655 133.415 ;
        RECT 93.280 133.370 93.570 133.415 ;
        RECT 96.060 133.370 96.350 133.415 ;
        RECT 97.920 133.370 98.210 133.415 ;
        RECT 81.365 133.230 88.020 133.370 ;
        RECT 81.365 133.185 81.655 133.230 ;
        RECT 50.530 133.030 50.850 133.090 ;
        RECT 46.940 132.890 50.850 133.030 ;
        RECT 44.090 132.830 44.410 132.890 ;
        RECT 44.565 132.845 44.855 132.890 ;
        RECT 50.530 132.830 50.850 132.890 ;
        RECT 80.445 133.030 80.735 133.075 ;
        RECT 83.190 133.030 83.510 133.090 ;
        RECT 80.445 132.890 83.510 133.030 ;
        RECT 87.880 133.030 88.020 133.230 ;
        RECT 93.280 133.230 98.210 133.370 ;
        RECT 100.300 133.370 100.440 133.570 ;
        RECT 100.670 133.510 100.990 133.770 ;
        RECT 102.050 133.710 102.370 133.770 ;
        RECT 104.825 133.710 105.115 133.755 ;
        RECT 102.050 133.570 105.115 133.710 ;
        RECT 102.050 133.510 102.370 133.570 ;
        RECT 104.825 133.525 105.115 133.570 ;
        RECT 109.500 133.370 109.640 133.850 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 100.300 133.230 109.640 133.370 ;
        RECT 93.280 133.185 93.570 133.230 ;
        RECT 96.060 133.185 96.350 133.230 ;
        RECT 97.920 133.185 98.210 133.230 ;
        RECT 94.690 133.030 95.010 133.090 ;
        RECT 87.880 132.890 95.010 133.030 ;
        RECT 80.445 132.845 80.735 132.890 ;
        RECT 83.190 132.830 83.510 132.890 ;
        RECT 94.690 132.830 95.010 132.890 ;
        RECT 98.845 133.030 99.135 133.075 ;
        RECT 99.750 133.030 100.070 133.090 ;
        RECT 98.845 132.890 100.070 133.030 ;
        RECT 98.845 132.845 99.135 132.890 ;
        RECT 99.750 132.830 100.070 132.890 ;
        RECT 101.130 132.830 101.450 133.090 ;
        RECT 103.430 132.830 103.750 133.090 ;
        RECT 104.810 132.830 105.130 133.090 ;
        RECT 109.885 133.030 110.175 133.075 ;
        RECT 110.330 133.030 110.650 133.090 ;
        RECT 109.885 132.890 110.650 133.030 ;
        RECT 109.885 132.845 110.175 132.890 ;
        RECT 110.330 132.830 110.650 132.890 ;
        RECT 111.250 132.830 111.570 133.090 ;
        RECT 14.580 132.210 127.740 132.690 ;
        RECT 28.910 131.810 29.230 132.070 ;
        RECT 30.750 132.055 31.070 132.070 ;
        RECT 30.535 131.825 31.070 132.055 ;
        RECT 30.750 131.810 31.070 131.825 ;
        RECT 33.970 132.010 34.290 132.070 ;
        RECT 78.605 132.010 78.895 132.055 ;
        RECT 79.970 132.010 80.290 132.070 ;
        RECT 33.970 131.870 40.180 132.010 ;
        RECT 33.970 131.810 34.290 131.870 ;
        RECT 40.040 131.730 40.180 131.870 ;
        RECT 78.605 131.870 80.290 132.010 ;
        RECT 78.605 131.825 78.895 131.870 ;
        RECT 79.970 131.810 80.290 131.870 ;
        RECT 89.645 132.010 89.935 132.055 ;
        RECT 90.550 132.010 90.870 132.070 ;
        RECT 89.645 131.870 90.870 132.010 ;
        RECT 89.645 131.825 89.935 131.870 ;
        RECT 90.550 131.810 90.870 131.870 ;
        RECT 109.870 131.810 110.190 132.070 ;
        RECT 34.400 131.670 34.690 131.715 ;
        RECT 37.180 131.670 37.470 131.715 ;
        RECT 39.040 131.670 39.330 131.715 ;
        RECT 34.400 131.530 39.330 131.670 ;
        RECT 34.400 131.485 34.690 131.530 ;
        RECT 37.180 131.485 37.470 131.530 ;
        RECT 39.040 131.485 39.330 131.530 ;
        RECT 39.950 131.670 40.270 131.730 ;
        RECT 69.865 131.670 70.155 131.715 ;
        RECT 100.210 131.670 100.530 131.730 ;
        RECT 39.950 131.530 100.530 131.670 ;
        RECT 39.950 131.470 40.270 131.530 ;
        RECT 69.865 131.485 70.155 131.530 ;
        RECT 100.210 131.470 100.530 131.530 ;
        RECT 102.510 131.670 102.830 131.730 ;
        RECT 118.150 131.670 118.470 131.730 ;
        RECT 102.510 131.530 118.470 131.670 ;
        RECT 102.510 131.470 102.830 131.530 ;
        RECT 118.150 131.470 118.470 131.530 ;
        RECT 21.105 131.330 21.395 131.375 ;
        RECT 22.010 131.330 22.330 131.390 ;
        RECT 21.105 131.190 22.330 131.330 ;
        RECT 21.105 131.145 21.395 131.190 ;
        RECT 22.010 131.130 22.330 131.190 ;
        RECT 36.270 131.330 36.590 131.390 ;
        RECT 36.270 131.190 37.420 131.330 ;
        RECT 36.270 131.130 36.590 131.190 ;
        RECT 28.450 130.990 28.770 131.050 ;
        RECT 29.845 130.990 30.135 131.035 ;
        RECT 28.450 130.850 30.135 130.990 ;
        RECT 28.450 130.790 28.770 130.850 ;
        RECT 29.845 130.805 30.135 130.850 ;
        RECT 34.400 130.990 34.690 131.035 ;
        RECT 37.280 130.990 37.420 131.190 ;
        RECT 37.650 131.130 37.970 131.390 ;
        RECT 64.790 131.330 65.110 131.390 ;
        RECT 66.645 131.330 66.935 131.375 ;
        RECT 69.390 131.330 69.710 131.390 ;
        RECT 64.790 131.190 69.710 131.330 ;
        RECT 64.790 131.130 65.110 131.190 ;
        RECT 66.645 131.145 66.935 131.190 ;
        RECT 69.390 131.130 69.710 131.190 ;
        RECT 73.545 131.330 73.835 131.375 ;
        RECT 73.990 131.330 74.310 131.390 ;
        RECT 73.545 131.190 74.310 131.330 ;
        RECT 73.545 131.145 73.835 131.190 ;
        RECT 73.990 131.130 74.310 131.190 ;
        RECT 39.505 130.990 39.795 131.035 ;
        RECT 70.785 130.990 71.075 131.035 ;
        RECT 72.610 130.990 72.930 131.050 ;
        RECT 74.465 130.990 74.755 131.035 ;
        RECT 79.525 130.990 79.815 131.035 ;
        RECT 34.400 130.850 36.935 130.990 ;
        RECT 37.280 130.850 42.480 130.990 ;
        RECT 34.400 130.805 34.690 130.850 ;
        RECT 22.025 130.650 22.315 130.695 ;
        RECT 23.390 130.650 23.710 130.710 ;
        RECT 22.025 130.510 23.710 130.650 ;
        RECT 22.025 130.465 22.315 130.510 ;
        RECT 23.390 130.450 23.710 130.510 ;
        RECT 32.540 130.650 32.830 130.695 ;
        RECT 33.970 130.650 34.290 130.710 ;
        RECT 36.720 130.695 36.935 130.850 ;
        RECT 39.505 130.805 39.795 130.850 ;
        RECT 35.800 130.650 36.090 130.695 ;
        RECT 32.540 130.510 36.090 130.650 ;
        RECT 32.540 130.465 32.830 130.510 ;
        RECT 33.970 130.450 34.290 130.510 ;
        RECT 35.800 130.465 36.090 130.510 ;
        RECT 36.720 130.650 37.010 130.695 ;
        RECT 38.580 130.650 38.870 130.695 ;
        RECT 36.720 130.510 38.870 130.650 ;
        RECT 36.720 130.465 37.010 130.510 ;
        RECT 38.580 130.465 38.870 130.510 ;
        RECT 21.565 130.310 21.855 130.355 ;
        RECT 22.470 130.310 22.790 130.370 ;
        RECT 21.565 130.170 22.790 130.310 ;
        RECT 21.565 130.125 21.855 130.170 ;
        RECT 22.470 130.110 22.790 130.170 ;
        RECT 22.930 130.310 23.250 130.370 ;
        RECT 42.340 130.355 42.480 130.850 ;
        RECT 70.785 130.850 74.755 130.990 ;
        RECT 70.785 130.805 71.075 130.850 ;
        RECT 72.610 130.790 72.930 130.850 ;
        RECT 74.465 130.805 74.755 130.850 ;
        RECT 75.000 130.850 79.815 130.990 ;
        RECT 48.705 130.650 48.995 130.695 ;
        RECT 49.150 130.650 49.470 130.710 ;
        RECT 48.705 130.510 49.470 130.650 ;
        RECT 48.705 130.465 48.995 130.510 ;
        RECT 49.150 130.450 49.470 130.510 ;
        RECT 64.330 130.650 64.650 130.710 ;
        RECT 65.710 130.650 66.030 130.710 ;
        RECT 67.565 130.650 67.855 130.695 ;
        RECT 64.330 130.510 67.855 130.650 ;
        RECT 64.330 130.450 64.650 130.510 ;
        RECT 65.710 130.450 66.030 130.510 ;
        RECT 67.565 130.465 67.855 130.510 ;
        RECT 68.010 130.650 68.330 130.710 ;
        RECT 75.000 130.650 75.140 130.850 ;
        RECT 79.525 130.805 79.815 130.850 ;
        RECT 79.970 130.790 80.290 131.050 ;
        RECT 88.250 130.990 88.570 131.050 ;
        RECT 89.185 130.990 89.475 131.035 ;
        RECT 91.010 130.990 91.330 131.050 ;
        RECT 88.250 130.850 91.330 130.990 ;
        RECT 88.250 130.790 88.570 130.850 ;
        RECT 89.185 130.805 89.475 130.850 ;
        RECT 91.010 130.790 91.330 130.850 ;
        RECT 98.370 130.990 98.690 131.050 ;
        RECT 100.225 130.990 100.515 131.035 ;
        RECT 98.370 130.850 100.515 130.990 ;
        RECT 98.370 130.790 98.690 130.850 ;
        RECT 100.225 130.805 100.515 130.850 ;
        RECT 110.790 130.790 111.110 131.050 ;
        RECT 111.725 130.990 112.015 131.035 ;
        RECT 112.170 130.990 112.490 131.050 ;
        RECT 111.725 130.850 112.490 130.990 ;
        RECT 111.725 130.805 112.015 130.850 ;
        RECT 112.170 130.790 112.490 130.850 ;
        RECT 68.010 130.510 75.140 130.650 ;
        RECT 68.010 130.450 68.330 130.510 ;
        RECT 75.000 130.370 75.140 130.510 ;
        RECT 23.865 130.310 24.155 130.355 ;
        RECT 22.930 130.170 24.155 130.310 ;
        RECT 22.930 130.110 23.250 130.170 ;
        RECT 23.865 130.125 24.155 130.170 ;
        RECT 42.265 130.310 42.555 130.355 ;
        RECT 42.710 130.310 43.030 130.370 ;
        RECT 42.265 130.170 43.030 130.310 ;
        RECT 42.265 130.125 42.555 130.170 ;
        RECT 42.710 130.110 43.030 130.170 ;
        RECT 66.170 130.310 66.490 130.370 ;
        RECT 67.105 130.310 67.395 130.355 ;
        RECT 66.170 130.170 67.395 130.310 ;
        RECT 66.170 130.110 66.490 130.170 ;
        RECT 67.105 130.125 67.395 130.170 ;
        RECT 69.405 130.310 69.695 130.355 ;
        RECT 70.310 130.310 70.630 130.370 ;
        RECT 69.405 130.170 70.630 130.310 ;
        RECT 69.405 130.125 69.695 130.170 ;
        RECT 70.310 130.110 70.630 130.170 ;
        RECT 71.690 130.110 72.010 130.370 ;
        RECT 74.910 130.110 75.230 130.370 ;
        RECT 14.580 129.490 127.740 129.970 ;
        RECT 17.655 129.290 17.945 129.335 ;
        RECT 23.390 129.290 23.710 129.350 ;
        RECT 17.655 129.150 27.760 129.290 ;
        RECT 17.655 129.105 17.945 129.150 ;
        RECT 23.390 129.090 23.710 129.150 ;
        RECT 19.660 128.950 19.950 128.995 ;
        RECT 21.090 128.950 21.410 129.010 ;
        RECT 22.920 128.950 23.210 128.995 ;
        RECT 19.660 128.810 23.210 128.950 ;
        RECT 19.660 128.765 19.950 128.810 ;
        RECT 21.090 128.750 21.410 128.810 ;
        RECT 22.920 128.765 23.210 128.810 ;
        RECT 23.840 128.950 24.130 128.995 ;
        RECT 25.700 128.950 25.990 128.995 ;
        RECT 23.840 128.810 25.990 128.950 ;
        RECT 27.620 128.950 27.760 129.150 ;
        RECT 33.970 129.090 34.290 129.350 ;
        RECT 37.650 129.290 37.970 129.350 ;
        RECT 38.585 129.290 38.875 129.335 ;
        RECT 37.650 129.150 38.875 129.290 ;
        RECT 37.650 129.090 37.970 129.150 ;
        RECT 38.585 129.105 38.875 129.150 ;
        RECT 41.805 129.290 42.095 129.335 ;
        RECT 43.630 129.290 43.950 129.350 ;
        RECT 41.805 129.150 43.950 129.290 ;
        RECT 41.805 129.105 42.095 129.150 ;
        RECT 43.630 129.090 43.950 129.150 ;
        RECT 44.105 129.290 44.395 129.335 ;
        RECT 45.010 129.290 45.330 129.350 ;
        RECT 44.105 129.150 45.330 129.290 ;
        RECT 44.105 129.105 44.395 129.150 ;
        RECT 45.010 129.090 45.330 129.150 ;
        RECT 49.165 129.290 49.455 129.335 ;
        RECT 49.610 129.290 49.930 129.350 ;
        RECT 49.165 129.150 49.930 129.290 ;
        RECT 49.165 129.105 49.455 129.150 ;
        RECT 49.610 129.090 49.930 129.150 ;
        RECT 55.590 129.290 55.910 129.350 ;
        RECT 56.065 129.290 56.355 129.335 ;
        RECT 55.590 129.150 56.355 129.290 ;
        RECT 55.590 129.090 55.910 129.150 ;
        RECT 56.065 129.105 56.355 129.150 ;
        RECT 56.510 129.090 56.830 129.350 ;
        RECT 65.035 129.290 65.325 129.335 ;
        RECT 66.170 129.290 66.490 129.350 ;
        RECT 65.035 129.150 66.490 129.290 ;
        RECT 65.035 129.105 65.325 129.150 ;
        RECT 66.170 129.090 66.490 129.150 ;
        RECT 77.760 129.150 81.580 129.290 ;
        RECT 42.710 128.950 43.030 129.010 ;
        RECT 46.865 128.950 47.155 128.995 ;
        RECT 63.870 128.950 64.190 129.010 ;
        RECT 27.620 128.810 40.180 128.950 ;
        RECT 23.840 128.765 24.130 128.810 ;
        RECT 25.700 128.765 25.990 128.810 ;
        RECT 21.520 128.610 21.810 128.655 ;
        RECT 23.840 128.610 24.055 128.765 ;
        RECT 21.520 128.470 24.055 128.610 ;
        RECT 26.625 128.610 26.915 128.655 ;
        RECT 29.830 128.610 30.150 128.670 ;
        RECT 26.625 128.470 30.150 128.610 ;
        RECT 21.520 128.425 21.810 128.470 ;
        RECT 26.625 128.425 26.915 128.470 ;
        RECT 29.830 128.410 30.150 128.470 ;
        RECT 30.290 128.610 30.610 128.670 ;
        RECT 33.525 128.610 33.815 128.655 ;
        RECT 30.290 128.470 33.815 128.610 ;
        RECT 30.290 128.410 30.610 128.470 ;
        RECT 33.525 128.425 33.815 128.470 ;
        RECT 39.490 128.410 39.810 128.670 ;
        RECT 40.040 128.655 40.180 128.810 ;
        RECT 42.710 128.810 64.190 128.950 ;
        RECT 42.710 128.750 43.030 128.810 ;
        RECT 46.865 128.765 47.155 128.810 ;
        RECT 63.870 128.750 64.190 128.810 ;
        RECT 67.040 128.950 67.330 128.995 ;
        RECT 68.470 128.950 68.790 129.010 ;
        RECT 70.300 128.950 70.590 128.995 ;
        RECT 67.040 128.810 70.590 128.950 ;
        RECT 67.040 128.765 67.330 128.810 ;
        RECT 68.470 128.750 68.790 128.810 ;
        RECT 70.300 128.765 70.590 128.810 ;
        RECT 71.220 128.950 71.510 128.995 ;
        RECT 73.080 128.950 73.370 128.995 ;
        RECT 71.220 128.810 73.370 128.950 ;
        RECT 71.220 128.765 71.510 128.810 ;
        RECT 73.080 128.765 73.370 128.810 ;
        RECT 39.965 128.425 40.255 128.655 ;
        RECT 40.885 128.610 41.175 128.655 ;
        RECT 43.185 128.610 43.475 128.655 ;
        RECT 45.930 128.610 46.250 128.670 ;
        RECT 48.245 128.610 48.535 128.655 ;
        RECT 68.010 128.610 68.330 128.670 ;
        RECT 40.885 128.470 68.330 128.610 ;
        RECT 40.885 128.425 41.175 128.470 ;
        RECT 43.185 128.425 43.475 128.470 ;
        RECT 45.930 128.410 46.250 128.470 ;
        RECT 48.245 128.425 48.535 128.470 ;
        RECT 68.010 128.410 68.330 128.470 ;
        RECT 68.900 128.610 69.190 128.655 ;
        RECT 71.220 128.610 71.435 128.765 ;
        RECT 68.900 128.470 71.435 128.610 ;
        RECT 68.900 128.425 69.190 128.470 ;
        RECT 72.150 128.410 72.470 128.670 ;
        RECT 74.910 128.610 75.230 128.670 ;
        RECT 77.760 128.655 77.900 129.150 ;
        RECT 78.605 128.950 78.895 128.995 ;
        RECT 80.430 128.950 80.750 129.010 ;
        RECT 78.605 128.810 80.750 128.950 ;
        RECT 81.440 128.950 81.580 129.150 ;
        RECT 83.190 129.090 83.510 129.350 ;
        RECT 88.250 129.090 88.570 129.350 ;
        RECT 89.645 129.105 89.935 129.335 ;
        RECT 81.440 128.810 84.340 128.950 ;
        RECT 78.605 128.765 78.895 128.810 ;
        RECT 80.430 128.750 80.750 128.810 ;
        RECT 84.200 128.655 84.340 128.810 ;
        RECT 84.660 128.810 85.720 128.950 ;
        RECT 75.385 128.610 75.675 128.655 ;
        RECT 77.685 128.610 77.975 128.655 ;
        RECT 80.905 128.610 81.195 128.655 ;
        RECT 74.910 128.470 77.975 128.610 ;
        RECT 74.910 128.410 75.230 128.470 ;
        RECT 75.385 128.425 75.675 128.470 ;
        RECT 77.685 128.425 77.975 128.470 ;
        RECT 79.140 128.470 81.195 128.610 ;
        RECT 23.850 128.270 24.170 128.330 ;
        RECT 24.785 128.270 25.075 128.315 ;
        RECT 23.850 128.130 25.075 128.270 ;
        RECT 23.850 128.070 24.170 128.130 ;
        RECT 24.785 128.085 25.075 128.130 ;
        RECT 42.265 128.085 42.555 128.315 ;
        RECT 42.710 128.270 43.030 128.330 ;
        RECT 47.325 128.270 47.615 128.315 ;
        RECT 42.710 128.130 47.615 128.270 ;
        RECT 21.520 127.930 21.810 127.975 ;
        RECT 24.300 127.930 24.590 127.975 ;
        RECT 26.160 127.930 26.450 127.975 ;
        RECT 21.520 127.790 26.450 127.930 ;
        RECT 21.520 127.745 21.810 127.790 ;
        RECT 24.300 127.745 24.590 127.790 ;
        RECT 26.160 127.745 26.450 127.790 ;
        RECT 22.470 127.590 22.790 127.650 ;
        RECT 42.340 127.590 42.480 128.085 ;
        RECT 42.710 128.070 43.030 128.130 ;
        RECT 47.325 128.085 47.615 128.130 ;
        RECT 54.670 128.270 54.990 128.330 ;
        RECT 55.145 128.270 55.435 128.315 ;
        RECT 54.670 128.130 55.435 128.270 ;
        RECT 54.670 128.070 54.990 128.130 ;
        RECT 55.145 128.085 55.435 128.130 ;
        RECT 63.870 128.270 64.190 128.330 ;
        RECT 74.005 128.270 74.295 128.315 ;
        RECT 63.870 128.130 74.295 128.270 ;
        RECT 63.870 128.070 64.190 128.130 ;
        RECT 74.005 128.085 74.295 128.130 ;
        RECT 74.465 128.085 74.755 128.315 ;
        RECT 76.765 128.270 77.055 128.315 ;
        RECT 78.590 128.270 78.910 128.330 ;
        RECT 79.140 128.270 79.280 128.470 ;
        RECT 80.905 128.425 81.195 128.470 ;
        RECT 84.125 128.425 84.415 128.655 ;
        RECT 76.765 128.130 79.280 128.270 ;
        RECT 76.765 128.085 77.055 128.130 ;
        RECT 68.900 127.930 69.190 127.975 ;
        RECT 71.680 127.930 71.970 127.975 ;
        RECT 73.540 127.930 73.830 127.975 ;
        RECT 68.900 127.790 73.830 127.930 ;
        RECT 74.540 127.930 74.680 128.085 ;
        RECT 78.590 128.070 78.910 128.130 ;
        RECT 79.985 128.085 80.275 128.315 ;
        RECT 79.050 127.930 79.370 127.990 ;
        RECT 74.540 127.790 79.370 127.930 ;
        RECT 80.060 127.930 80.200 128.085 ;
        RECT 80.430 128.070 80.750 128.330 ;
        RECT 80.980 128.270 81.120 128.425 ;
        RECT 84.660 128.270 84.800 128.810 ;
        RECT 85.045 128.425 85.335 128.655 ;
        RECT 80.980 128.130 84.800 128.270 ;
        RECT 85.120 127.930 85.260 128.425 ;
        RECT 85.580 128.270 85.720 128.810 ;
        RECT 87.345 128.610 87.635 128.655 ;
        RECT 89.720 128.610 89.860 129.105 ;
        RECT 95.150 129.090 95.470 129.350 ;
        RECT 98.370 129.290 98.690 129.350 ;
        RECT 102.065 129.290 102.355 129.335 ;
        RECT 98.370 129.150 102.355 129.290 ;
        RECT 98.370 129.090 98.690 129.150 ;
        RECT 102.065 129.105 102.355 129.150 ;
        RECT 104.810 129.090 105.130 129.350 ;
        RECT 106.190 129.290 106.510 129.350 ;
        RECT 107.125 129.290 107.415 129.335 ;
        RECT 106.190 129.150 107.415 129.290 ;
        RECT 106.190 129.090 106.510 129.150 ;
        RECT 107.125 129.105 107.415 129.150 ;
        RECT 111.250 129.090 111.570 129.350 ;
        RECT 95.610 128.750 95.930 129.010 ;
        RECT 105.820 128.810 108.260 128.950 ;
        RECT 87.345 128.470 89.860 128.610 ;
        RECT 91.485 128.610 91.775 128.655 ;
        RECT 93.770 128.610 94.090 128.670 ;
        RECT 94.245 128.610 94.535 128.655 ;
        RECT 91.485 128.470 93.540 128.610 ;
        RECT 87.345 128.425 87.635 128.470 ;
        RECT 91.485 128.425 91.775 128.470 ;
        RECT 91.945 128.270 92.235 128.315 ;
        RECT 85.580 128.130 92.235 128.270 ;
        RECT 91.945 128.085 92.235 128.130 ;
        RECT 92.405 128.085 92.695 128.315 ;
        RECT 93.400 128.270 93.540 128.470 ;
        RECT 93.770 128.470 94.535 128.610 ;
        RECT 93.770 128.410 94.090 128.470 ;
        RECT 94.245 128.425 94.535 128.470 ;
        RECT 100.210 128.610 100.530 128.670 ;
        RECT 105.820 128.655 105.960 128.810 ;
        RECT 105.745 128.610 106.035 128.655 ;
        RECT 100.210 128.470 106.035 128.610 ;
        RECT 100.210 128.410 100.530 128.470 ;
        RECT 105.745 128.425 106.035 128.470 ;
        RECT 106.190 128.410 106.510 128.670 ;
        RECT 108.120 128.655 108.260 128.810 ;
        RECT 108.045 128.610 108.335 128.655 ;
        RECT 110.345 128.610 110.635 128.655 ;
        RECT 110.790 128.610 111.110 128.670 ;
        RECT 112.645 128.610 112.935 128.655 ;
        RECT 108.045 128.470 112.935 128.610 ;
        RECT 108.045 128.425 108.335 128.470 ;
        RECT 110.345 128.425 110.635 128.470 ;
        RECT 110.790 128.410 111.110 128.470 ;
        RECT 112.645 128.425 112.935 128.470 ;
        RECT 113.090 128.410 113.410 128.670 ;
        RECT 118.150 128.410 118.470 128.670 ;
        RECT 119.545 128.425 119.835 128.655 ;
        RECT 98.830 128.270 99.150 128.330 ;
        RECT 105.270 128.270 105.590 128.330 ;
        RECT 108.965 128.270 109.255 128.315 ;
        RECT 93.400 128.130 109.255 128.270 ;
        RECT 91.470 127.930 91.790 127.990 ;
        RECT 80.060 127.790 84.800 127.930 ;
        RECT 85.120 127.790 91.790 127.930 ;
        RECT 68.900 127.745 69.190 127.790 ;
        RECT 71.680 127.745 71.970 127.790 ;
        RECT 73.540 127.745 73.830 127.790 ;
        RECT 79.050 127.730 79.370 127.790 ;
        RECT 84.660 127.650 84.800 127.790 ;
        RECT 91.470 127.730 91.790 127.790 ;
        RECT 22.470 127.450 42.480 127.590 ;
        RECT 57.890 127.590 58.210 127.650 ;
        RECT 58.365 127.590 58.655 127.635 ;
        RECT 57.890 127.450 58.655 127.590 ;
        RECT 22.470 127.390 22.790 127.450 ;
        RECT 57.890 127.390 58.210 127.450 ;
        RECT 58.365 127.405 58.655 127.450 ;
        RECT 76.305 127.590 76.595 127.635 ;
        RECT 81.810 127.590 82.130 127.650 ;
        RECT 76.305 127.450 82.130 127.590 ;
        RECT 76.305 127.405 76.595 127.450 ;
        RECT 81.810 127.390 82.130 127.450 ;
        RECT 82.745 127.590 83.035 127.635 ;
        RECT 83.650 127.590 83.970 127.650 ;
        RECT 82.745 127.450 83.970 127.590 ;
        RECT 82.745 127.405 83.035 127.450 ;
        RECT 83.650 127.390 83.970 127.450 ;
        RECT 84.570 127.590 84.890 127.650 ;
        RECT 92.480 127.590 92.620 128.085 ;
        RECT 98.830 128.070 99.150 128.130 ;
        RECT 105.270 128.070 105.590 128.130 ;
        RECT 108.965 128.085 109.255 128.130 ;
        RECT 109.410 128.070 109.730 128.330 ;
        RECT 114.930 128.270 115.250 128.330 ;
        RECT 119.620 128.270 119.760 128.425 ;
        RECT 114.930 128.130 119.760 128.270 ;
        RECT 114.930 128.070 115.250 128.130 ;
        RECT 102.970 127.930 103.290 127.990 ;
        RECT 111.725 127.930 112.015 127.975 ;
        RECT 102.970 127.790 112.015 127.930 ;
        RECT 102.970 127.730 103.290 127.790 ;
        RECT 111.725 127.745 112.015 127.790 ;
        RECT 84.570 127.450 92.620 127.590 ;
        RECT 84.570 127.390 84.890 127.450 ;
        RECT 118.610 127.390 118.930 127.650 ;
        RECT 120.450 127.390 120.770 127.650 ;
        RECT 14.580 126.770 127.740 127.250 ;
        RECT 23.850 126.370 24.170 126.630 ;
        RECT 71.245 126.570 71.535 126.615 ;
        RECT 72.150 126.570 72.470 126.630 ;
        RECT 78.590 126.615 78.910 126.630 ;
        RECT 71.245 126.430 72.470 126.570 ;
        RECT 71.245 126.385 71.535 126.430 ;
        RECT 72.150 126.370 72.470 126.430 ;
        RECT 78.375 126.385 78.910 126.615 ;
        RECT 78.590 126.370 78.910 126.385 ;
        RECT 79.050 126.570 79.370 126.630 ;
        RECT 80.430 126.570 80.750 126.630 ;
        RECT 98.830 126.615 99.150 126.630 ;
        RECT 79.050 126.430 80.750 126.570 ;
        RECT 79.050 126.370 79.370 126.430 ;
        RECT 80.430 126.370 80.750 126.430 ;
        RECT 98.615 126.385 99.150 126.615 ;
        RECT 98.830 126.370 99.150 126.385 ;
        RECT 114.930 126.370 115.250 126.630 ;
        RECT 55.590 126.230 55.910 126.290 ;
        RECT 82.240 126.230 82.530 126.275 ;
        RECT 85.020 126.230 85.310 126.275 ;
        RECT 86.880 126.230 87.170 126.275 ;
        RECT 55.590 126.090 60.880 126.230 ;
        RECT 55.590 126.030 55.910 126.090 ;
        RECT 19.710 125.890 20.030 125.950 ;
        RECT 30.290 125.890 30.610 125.950 ;
        RECT 19.710 125.750 30.610 125.890 ;
        RECT 19.710 125.690 20.030 125.750 ;
        RECT 21.090 125.550 21.410 125.610 ;
        RECT 22.100 125.595 22.240 125.750 ;
        RECT 30.290 125.690 30.610 125.750 ;
        RECT 35.810 125.890 36.130 125.950 ;
        RECT 42.725 125.890 43.015 125.935 ;
        RECT 54.670 125.890 54.990 125.950 ;
        RECT 59.745 125.890 60.035 125.935 ;
        RECT 35.810 125.750 43.015 125.890 ;
        RECT 35.810 125.690 36.130 125.750 ;
        RECT 42.725 125.705 43.015 125.750 ;
        RECT 43.720 125.750 46.160 125.890 ;
        RECT 21.565 125.550 21.855 125.595 ;
        RECT 21.090 125.410 21.855 125.550 ;
        RECT 21.090 125.350 21.410 125.410 ;
        RECT 21.565 125.365 21.855 125.410 ;
        RECT 22.025 125.365 22.315 125.595 ;
        RECT 22.930 125.350 23.250 125.610 ;
        RECT 36.730 125.350 37.050 125.610 ;
        RECT 37.665 125.365 37.955 125.595 ;
        RECT 38.110 125.550 38.430 125.610 ;
        RECT 38.585 125.550 38.875 125.595 ;
        RECT 38.110 125.410 38.875 125.550 ;
        RECT 37.740 125.210 37.880 125.365 ;
        RECT 38.110 125.350 38.430 125.410 ;
        RECT 38.585 125.365 38.875 125.410 ;
        RECT 40.410 125.350 40.730 125.610 ;
        RECT 41.345 125.365 41.635 125.595 ;
        RECT 39.950 125.210 40.270 125.270 ;
        RECT 37.740 125.070 40.270 125.210 ;
        RECT 41.420 125.210 41.560 125.365 ;
        RECT 42.250 125.350 42.570 125.610 ;
        RECT 43.720 125.595 43.860 125.750 ;
        RECT 46.020 125.610 46.160 125.750 ;
        RECT 54.670 125.750 60.035 125.890 ;
        RECT 60.740 125.890 60.880 126.090 ;
        RECT 82.240 126.090 87.170 126.230 ;
        RECT 82.240 126.045 82.530 126.090 ;
        RECT 85.020 126.045 85.310 126.090 ;
        RECT 86.880 126.045 87.170 126.090 ;
        RECT 90.110 126.230 90.400 126.275 ;
        RECT 91.970 126.230 92.260 126.275 ;
        RECT 94.750 126.230 95.040 126.275 ;
        RECT 90.110 126.090 95.040 126.230 ;
        RECT 90.110 126.045 90.400 126.090 ;
        RECT 91.970 126.045 92.260 126.090 ;
        RECT 94.750 126.045 95.040 126.090 ;
        RECT 119.500 126.230 119.790 126.275 ;
        RECT 122.280 126.230 122.570 126.275 ;
        RECT 124.140 126.230 124.430 126.275 ;
        RECT 119.500 126.090 124.430 126.230 ;
        RECT 119.500 126.045 119.790 126.090 ;
        RECT 122.280 126.045 122.570 126.090 ;
        RECT 124.140 126.045 124.430 126.090 ;
        RECT 74.465 125.890 74.755 125.935 ;
        RECT 79.510 125.890 79.830 125.950 ;
        RECT 84.570 125.890 84.890 125.950 ;
        RECT 60.740 125.750 61.340 125.890 ;
        RECT 54.670 125.690 54.990 125.750 ;
        RECT 59.745 125.705 60.035 125.750 ;
        RECT 43.645 125.550 43.935 125.595 ;
        RECT 42.800 125.410 43.935 125.550 ;
        RECT 42.800 125.210 42.940 125.410 ;
        RECT 43.645 125.365 43.935 125.410 ;
        RECT 44.550 125.350 44.870 125.610 ;
        RECT 45.930 125.350 46.250 125.610 ;
        RECT 46.390 125.350 46.710 125.610 ;
        RECT 57.890 125.350 58.210 125.610 ;
        RECT 60.650 125.350 60.970 125.610 ;
        RECT 61.200 125.595 61.340 125.750 ;
        RECT 74.465 125.750 84.890 125.890 ;
        RECT 74.465 125.705 74.755 125.750 ;
        RECT 79.510 125.690 79.830 125.750 ;
        RECT 84.570 125.690 84.890 125.750 ;
        RECT 88.250 125.890 88.570 125.950 ;
        RECT 91.485 125.890 91.775 125.935 ;
        RECT 98.370 125.890 98.690 125.950 ;
        RECT 88.250 125.750 91.775 125.890 ;
        RECT 88.250 125.690 88.570 125.750 ;
        RECT 91.485 125.705 91.775 125.750 ;
        RECT 92.020 125.750 98.690 125.890 ;
        RECT 61.125 125.365 61.415 125.595 ;
        RECT 68.470 125.550 68.790 125.610 ;
        RECT 68.945 125.550 69.235 125.595 ;
        RECT 68.470 125.410 69.235 125.550 ;
        RECT 68.470 125.350 68.790 125.410 ;
        RECT 68.945 125.365 69.235 125.410 ;
        RECT 69.405 125.550 69.695 125.595 ;
        RECT 69.850 125.550 70.170 125.610 ;
        RECT 69.405 125.410 70.170 125.550 ;
        RECT 69.405 125.365 69.695 125.410 ;
        RECT 69.850 125.350 70.170 125.410 ;
        RECT 70.310 125.350 70.630 125.610 ;
        RECT 71.690 125.550 72.010 125.610 ;
        RECT 73.085 125.550 73.375 125.595 ;
        RECT 71.090 125.410 73.375 125.550 ;
        RECT 41.420 125.070 42.940 125.210 ;
        RECT 43.170 125.210 43.490 125.270 ;
        RECT 45.025 125.210 45.315 125.255 ;
        RECT 43.170 125.070 45.315 125.210 ;
        RECT 39.950 125.010 40.270 125.070 ;
        RECT 43.170 125.010 43.490 125.070 ;
        RECT 45.025 125.025 45.315 125.070 ;
        RECT 49.165 125.210 49.455 125.255 ;
        RECT 71.090 125.210 71.230 125.410 ;
        RECT 71.690 125.350 72.010 125.410 ;
        RECT 73.085 125.365 73.375 125.410 ;
        RECT 82.240 125.550 82.530 125.595 ;
        RECT 82.240 125.410 84.775 125.550 ;
        RECT 82.240 125.365 82.530 125.410 ;
        RECT 49.165 125.070 71.230 125.210 ;
        RECT 80.380 125.210 80.670 125.255 ;
        RECT 82.730 125.210 83.050 125.270 ;
        RECT 84.560 125.255 84.775 125.410 ;
        RECT 85.490 125.350 85.810 125.610 ;
        RECT 87.345 125.550 87.635 125.595 ;
        RECT 89.645 125.550 89.935 125.595 ;
        RECT 92.020 125.550 92.160 125.750 ;
        RECT 98.370 125.690 98.690 125.750 ;
        RECT 112.185 125.890 112.475 125.935 ;
        RECT 113.550 125.890 113.870 125.950 ;
        RECT 112.185 125.750 113.870 125.890 ;
        RECT 112.185 125.705 112.475 125.750 ;
        RECT 113.550 125.690 113.870 125.750 ;
        RECT 120.450 125.890 120.770 125.950 ;
        RECT 122.765 125.890 123.055 125.935 ;
        RECT 120.450 125.750 123.055 125.890 ;
        RECT 120.450 125.690 120.770 125.750 ;
        RECT 122.765 125.705 123.055 125.750 ;
        RECT 94.750 125.550 95.040 125.595 ;
        RECT 87.345 125.410 92.160 125.550 ;
        RECT 92.505 125.410 95.040 125.550 ;
        RECT 87.345 125.365 87.635 125.410 ;
        RECT 89.645 125.365 89.935 125.410 ;
        RECT 92.505 125.255 92.720 125.410 ;
        RECT 94.750 125.365 95.040 125.410 ;
        RECT 99.290 125.350 99.610 125.610 ;
        RECT 100.210 125.350 100.530 125.610 ;
        RECT 101.130 125.350 101.450 125.610 ;
        RECT 105.270 125.550 105.590 125.610 ;
        RECT 112.645 125.550 112.935 125.595 ;
        RECT 105.270 125.410 112.935 125.550 ;
        RECT 105.270 125.350 105.590 125.410 ;
        RECT 112.645 125.365 112.935 125.410 ;
        RECT 119.500 125.550 119.790 125.595 ;
        RECT 119.500 125.410 122.035 125.550 ;
        RECT 119.500 125.365 119.790 125.410 ;
        RECT 83.640 125.210 83.930 125.255 ;
        RECT 80.380 125.070 83.930 125.210 ;
        RECT 49.165 125.025 49.455 125.070 ;
        RECT 80.380 125.025 80.670 125.070 ;
        RECT 82.730 125.010 83.050 125.070 ;
        RECT 83.640 125.025 83.930 125.070 ;
        RECT 84.560 125.210 84.850 125.255 ;
        RECT 86.420 125.210 86.710 125.255 ;
        RECT 84.560 125.070 86.710 125.210 ;
        RECT 84.560 125.025 84.850 125.070 ;
        RECT 86.420 125.025 86.710 125.070 ;
        RECT 90.570 125.210 90.860 125.255 ;
        RECT 92.430 125.210 92.720 125.255 ;
        RECT 90.570 125.070 92.720 125.210 ;
        RECT 90.570 125.025 90.860 125.070 ;
        RECT 92.430 125.025 92.720 125.070 ;
        RECT 93.310 125.255 93.630 125.270 ;
        RECT 93.310 125.210 93.640 125.255 ;
        RECT 96.610 125.210 96.900 125.255 ;
        RECT 93.310 125.070 96.900 125.210 ;
        RECT 93.310 125.025 93.640 125.070 ;
        RECT 96.610 125.025 96.900 125.070 ;
        RECT 117.640 125.210 117.930 125.255 ;
        RECT 118.610 125.210 118.930 125.270 ;
        RECT 121.820 125.255 122.035 125.410 ;
        RECT 124.590 125.350 124.910 125.610 ;
        RECT 120.900 125.210 121.190 125.255 ;
        RECT 117.640 125.070 121.190 125.210 ;
        RECT 117.640 125.025 117.930 125.070 ;
        RECT 93.310 125.010 93.630 125.025 ;
        RECT 118.610 125.010 118.930 125.070 ;
        RECT 120.900 125.025 121.190 125.070 ;
        RECT 121.820 125.210 122.110 125.255 ;
        RECT 123.680 125.210 123.970 125.255 ;
        RECT 121.820 125.070 123.970 125.210 ;
        RECT 121.820 125.025 122.110 125.070 ;
        RECT 123.680 125.025 123.970 125.070 ;
        RECT 45.930 124.870 46.250 124.930 ;
        RECT 47.785 124.870 48.075 124.915 ;
        RECT 45.930 124.730 48.075 124.870 ;
        RECT 45.930 124.670 46.250 124.730 ;
        RECT 47.785 124.685 48.075 124.730 ;
        RECT 58.825 124.870 59.115 124.915 ;
        RECT 60.190 124.870 60.510 124.930 ;
        RECT 58.825 124.730 60.510 124.870 ;
        RECT 58.825 124.685 59.115 124.730 ;
        RECT 60.190 124.670 60.510 124.730 ;
        RECT 62.965 124.870 63.255 124.915 ;
        RECT 69.850 124.870 70.170 124.930 ;
        RECT 62.965 124.730 70.170 124.870 ;
        RECT 62.965 124.685 63.255 124.730 ;
        RECT 69.850 124.670 70.170 124.730 ;
        RECT 113.090 124.870 113.410 124.930 ;
        RECT 115.635 124.870 115.925 124.915 ;
        RECT 113.090 124.730 115.925 124.870 ;
        RECT 113.090 124.670 113.410 124.730 ;
        RECT 115.635 124.685 115.925 124.730 ;
        RECT 14.580 124.050 127.740 124.530 ;
        RECT 22.470 123.850 22.790 123.910 ;
        RECT 23.390 123.850 23.710 123.910 ;
        RECT 24.325 123.850 24.615 123.895 ;
        RECT 22.470 123.650 22.930 123.850 ;
        RECT 23.390 123.710 24.615 123.850 ;
        RECT 23.390 123.650 23.710 123.710 ;
        RECT 24.325 123.665 24.615 123.710 ;
        RECT 24.785 123.850 25.075 123.895 ;
        RECT 42.710 123.850 43.030 123.910 ;
        RECT 24.785 123.710 43.030 123.850 ;
        RECT 24.785 123.665 25.075 123.710 ;
        RECT 22.790 123.510 22.930 123.650 ;
        RECT 24.860 123.510 25.000 123.665 ;
        RECT 42.710 123.650 43.030 123.710 ;
        RECT 53.075 123.850 53.365 123.895 ;
        RECT 55.590 123.850 55.910 123.910 ;
        RECT 53.075 123.710 55.910 123.850 ;
        RECT 53.075 123.665 53.365 123.710 ;
        RECT 55.590 123.650 55.910 123.710 ;
        RECT 60.650 123.850 60.970 123.910 ;
        RECT 65.725 123.850 66.015 123.895 ;
        RECT 60.650 123.710 66.015 123.850 ;
        RECT 60.650 123.650 60.970 123.710 ;
        RECT 65.725 123.665 66.015 123.710 ;
        RECT 82.285 123.850 82.575 123.895 ;
        RECT 82.730 123.850 83.050 123.910 ;
        RECT 82.285 123.710 83.050 123.850 ;
        RECT 82.285 123.665 82.575 123.710 ;
        RECT 82.730 123.650 83.050 123.710 ;
        RECT 84.585 123.850 84.875 123.895 ;
        RECT 85.490 123.850 85.810 123.910 ;
        RECT 84.585 123.710 85.810 123.850 ;
        RECT 84.585 123.665 84.875 123.710 ;
        RECT 85.490 123.650 85.810 123.710 ;
        RECT 93.310 123.650 93.630 123.910 ;
        RECT 22.790 123.370 25.000 123.510 ;
        RECT 55.080 123.510 55.370 123.555 ;
        RECT 57.430 123.510 57.750 123.570 ;
        RECT 58.340 123.510 58.630 123.555 ;
        RECT 55.080 123.370 58.630 123.510 ;
        RECT 55.080 123.325 55.370 123.370 ;
        RECT 57.430 123.310 57.750 123.370 ;
        RECT 58.340 123.325 58.630 123.370 ;
        RECT 59.260 123.510 59.550 123.555 ;
        RECT 61.120 123.510 61.410 123.555 ;
        RECT 59.260 123.370 61.410 123.510 ;
        RECT 59.260 123.325 59.550 123.370 ;
        RECT 61.120 123.325 61.410 123.370 ;
        RECT 111.725 123.510 112.015 123.555 ;
        RECT 113.090 123.510 113.410 123.570 ;
        RECT 111.725 123.370 113.410 123.510 ;
        RECT 111.725 123.325 112.015 123.370 ;
        RECT 34.890 122.970 35.210 123.230 ;
        RECT 56.940 123.170 57.230 123.215 ;
        RECT 59.260 123.170 59.475 123.325 ;
        RECT 113.090 123.310 113.410 123.370 ;
        RECT 117.640 123.510 117.930 123.555 ;
        RECT 119.070 123.510 119.390 123.570 ;
        RECT 120.900 123.510 121.190 123.555 ;
        RECT 117.640 123.370 121.190 123.510 ;
        RECT 117.640 123.325 117.930 123.370 ;
        RECT 119.070 123.310 119.390 123.370 ;
        RECT 120.900 123.325 121.190 123.370 ;
        RECT 121.820 123.510 122.110 123.555 ;
        RECT 123.680 123.510 123.970 123.555 ;
        RECT 121.820 123.370 123.970 123.510 ;
        RECT 121.820 123.325 122.110 123.370 ;
        RECT 123.680 123.325 123.970 123.370 ;
        RECT 56.940 123.030 59.475 123.170 ;
        RECT 56.940 122.985 57.230 123.030 ;
        RECT 60.190 122.970 60.510 123.230 ;
        RECT 62.045 123.170 62.335 123.215 ;
        RECT 63.870 123.170 64.190 123.230 ;
        RECT 62.045 123.030 64.190 123.170 ;
        RECT 62.045 122.985 62.335 123.030 ;
        RECT 63.870 122.970 64.190 123.030 ;
        RECT 64.330 123.170 64.650 123.230 ;
        RECT 65.265 123.170 65.555 123.215 ;
        RECT 64.330 123.030 65.555 123.170 ;
        RECT 64.330 122.970 64.650 123.030 ;
        RECT 65.265 122.985 65.555 123.030 ;
        RECT 73.070 123.170 73.390 123.230 ;
        RECT 82.745 123.170 83.035 123.215 ;
        RECT 83.190 123.170 83.510 123.230 ;
        RECT 73.070 123.030 83.510 123.170 ;
        RECT 73.070 122.970 73.390 123.030 ;
        RECT 82.745 122.985 83.035 123.030 ;
        RECT 83.190 122.970 83.510 123.030 ;
        RECT 83.650 122.970 83.970 123.230 ;
        RECT 91.010 123.170 91.330 123.230 ;
        RECT 92.865 123.170 93.155 123.215 ;
        RECT 100.210 123.170 100.530 123.230 ;
        RECT 91.010 123.030 100.530 123.170 ;
        RECT 91.010 122.970 91.330 123.030 ;
        RECT 92.865 122.985 93.155 123.030 ;
        RECT 100.210 122.970 100.530 123.030 ;
        RECT 112.185 123.170 112.475 123.215 ;
        RECT 112.630 123.170 112.950 123.230 ;
        RECT 115.635 123.170 115.925 123.215 ;
        RECT 112.185 123.030 115.925 123.170 ;
        RECT 112.185 122.985 112.475 123.030 ;
        RECT 112.630 122.970 112.950 123.030 ;
        RECT 115.635 122.985 115.925 123.030 ;
        RECT 119.500 123.170 119.790 123.215 ;
        RECT 121.820 123.170 122.035 123.325 ;
        RECT 119.500 123.030 122.035 123.170 ;
        RECT 119.500 122.985 119.790 123.030 ;
        RECT 124.590 122.970 124.910 123.230 ;
        RECT 22.010 122.830 22.330 122.890 ;
        RECT 23.405 122.830 23.695 122.875 ;
        RECT 33.525 122.830 33.815 122.875 ;
        RECT 22.010 122.690 33.815 122.830 ;
        RECT 22.010 122.630 22.330 122.690 ;
        RECT 23.405 122.645 23.695 122.690 ;
        RECT 33.525 122.645 33.815 122.690 ;
        RECT 34.445 122.830 34.735 122.875 ;
        RECT 36.730 122.830 37.050 122.890 ;
        RECT 41.790 122.830 42.110 122.890 ;
        RECT 34.445 122.690 42.110 122.830 ;
        RECT 34.445 122.645 34.735 122.690 ;
        RECT 33.600 122.490 33.740 122.645 ;
        RECT 36.730 122.630 37.050 122.690 ;
        RECT 41.790 122.630 42.110 122.690 ;
        RECT 64.790 122.630 65.110 122.890 ;
        RECT 105.270 122.830 105.590 122.890 ;
        RECT 110.805 122.830 111.095 122.875 ;
        RECT 113.550 122.830 113.870 122.890 ;
        RECT 105.270 122.690 113.870 122.830 ;
        RECT 105.270 122.630 105.590 122.690 ;
        RECT 110.805 122.645 111.095 122.690 ;
        RECT 113.550 122.630 113.870 122.690 ;
        RECT 121.370 122.830 121.690 122.890 ;
        RECT 122.765 122.830 123.055 122.875 ;
        RECT 121.370 122.690 123.055 122.830 ;
        RECT 121.370 122.630 121.690 122.690 ;
        RECT 122.765 122.645 123.055 122.690 ;
        RECT 43.630 122.490 43.950 122.550 ;
        RECT 45.930 122.490 46.250 122.550 ;
        RECT 46.850 122.490 47.170 122.550 ;
        RECT 33.600 122.350 47.170 122.490 ;
        RECT 43.630 122.290 43.950 122.350 ;
        RECT 45.930 122.290 46.250 122.350 ;
        RECT 46.850 122.290 47.170 122.350 ;
        RECT 56.940 122.490 57.230 122.535 ;
        RECT 59.720 122.490 60.010 122.535 ;
        RECT 61.580 122.490 61.870 122.535 ;
        RECT 56.940 122.350 61.870 122.490 ;
        RECT 56.940 122.305 57.230 122.350 ;
        RECT 59.720 122.305 60.010 122.350 ;
        RECT 61.580 122.305 61.870 122.350 ;
        RECT 119.500 122.490 119.790 122.535 ;
        RECT 122.280 122.490 122.570 122.535 ;
        RECT 124.140 122.490 124.430 122.535 ;
        RECT 119.500 122.350 124.430 122.490 ;
        RECT 119.500 122.305 119.790 122.350 ;
        RECT 122.280 122.305 122.570 122.350 ;
        RECT 124.140 122.305 124.430 122.350 ;
        RECT 26.610 121.950 26.930 122.210 ;
        RECT 36.730 121.950 37.050 122.210 ;
        RECT 67.565 122.150 67.855 122.195 ;
        RECT 68.010 122.150 68.330 122.210 ;
        RECT 67.565 122.010 68.330 122.150 ;
        RECT 67.565 121.965 67.855 122.010 ;
        RECT 68.010 121.950 68.330 122.010 ;
        RECT 114.025 122.150 114.315 122.195 ;
        RECT 120.450 122.150 120.770 122.210 ;
        RECT 114.025 122.010 120.770 122.150 ;
        RECT 114.025 121.965 114.315 122.010 ;
        RECT 120.450 121.950 120.770 122.010 ;
        RECT 14.580 121.330 127.740 121.810 ;
        RECT 30.535 121.130 30.825 121.175 ;
        RECT 34.890 121.130 35.210 121.190 ;
        RECT 30.535 120.990 35.210 121.130 ;
        RECT 30.535 120.945 30.825 120.990 ;
        RECT 34.890 120.930 35.210 120.990 ;
        RECT 57.430 120.930 57.750 121.190 ;
        RECT 59.515 121.130 59.805 121.175 ;
        RECT 60.650 121.130 60.970 121.190 ;
        RECT 59.515 120.990 60.970 121.130 ;
        RECT 59.515 120.945 59.805 120.990 ;
        RECT 60.650 120.930 60.970 120.990 ;
        RECT 119.070 120.930 119.390 121.190 ;
        RECT 121.370 120.930 121.690 121.190 ;
        RECT 22.010 120.790 22.330 120.850 ;
        RECT 34.400 120.790 34.690 120.835 ;
        RECT 37.180 120.790 37.470 120.835 ;
        RECT 39.040 120.790 39.330 120.835 ;
        RECT 63.380 120.790 63.670 120.835 ;
        RECT 66.160 120.790 66.450 120.835 ;
        RECT 68.020 120.790 68.310 120.835 ;
        RECT 22.010 120.650 23.160 120.790 ;
        RECT 22.010 120.590 22.330 120.650 ;
        RECT 22.470 120.250 22.790 120.510 ;
        RECT 23.020 120.495 23.160 120.650 ;
        RECT 34.400 120.650 39.330 120.790 ;
        RECT 34.400 120.605 34.690 120.650 ;
        RECT 37.180 120.605 37.470 120.650 ;
        RECT 39.040 120.605 39.330 120.650 ;
        RECT 42.800 120.650 47.540 120.790 ;
        RECT 22.945 120.265 23.235 120.495 ;
        RECT 35.810 120.450 36.130 120.510 ;
        RECT 42.800 120.450 42.940 120.650 ;
        RECT 30.840 120.310 42.940 120.450 ;
        RECT 43.185 120.450 43.475 120.495 ;
        RECT 43.630 120.450 43.950 120.510 ;
        RECT 43.185 120.310 43.950 120.450 ;
        RECT 26.610 120.110 26.930 120.170 ;
        RECT 27.085 120.110 27.375 120.155 ;
        RECT 26.610 119.970 27.375 120.110 ;
        RECT 26.610 119.910 26.930 119.970 ;
        RECT 27.085 119.925 27.375 119.970 ;
        RECT 30.840 119.830 30.980 120.310 ;
        RECT 35.810 120.250 36.130 120.310 ;
        RECT 43.185 120.265 43.475 120.310 ;
        RECT 43.630 120.250 43.950 120.310 ;
        RECT 46.390 120.250 46.710 120.510 ;
        RECT 46.850 120.250 47.170 120.510 ;
        RECT 47.400 120.495 47.540 120.650 ;
        RECT 63.380 120.650 68.310 120.790 ;
        RECT 63.380 120.605 63.670 120.650 ;
        RECT 66.160 120.605 66.450 120.650 ;
        RECT 68.020 120.605 68.310 120.650 ;
        RECT 68.945 120.605 69.235 120.835 ;
        RECT 113.060 120.790 113.350 120.835 ;
        RECT 115.840 120.790 116.130 120.835 ;
        RECT 117.700 120.790 117.990 120.835 ;
        RECT 113.060 120.650 117.990 120.790 ;
        RECT 113.060 120.605 113.350 120.650 ;
        RECT 115.840 120.605 116.130 120.650 ;
        RECT 117.700 120.605 117.990 120.650 ;
        RECT 47.325 120.265 47.615 120.495 ;
        RECT 66.645 120.450 66.935 120.495 ;
        RECT 69.020 120.450 69.160 120.605 ;
        RECT 66.645 120.310 69.160 120.450 ;
        RECT 77.685 120.450 77.975 120.495 ;
        RECT 79.510 120.450 79.830 120.510 ;
        RECT 83.650 120.450 83.970 120.510 ;
        RECT 93.785 120.450 94.075 120.495 ;
        RECT 97.925 120.450 98.215 120.495 ;
        RECT 105.270 120.450 105.590 120.510 ;
        RECT 109.410 120.495 109.730 120.510 ;
        RECT 77.685 120.310 105.590 120.450 ;
        RECT 66.645 120.265 66.935 120.310 ;
        RECT 77.685 120.265 77.975 120.310 ;
        RECT 79.510 120.250 79.830 120.310 ;
        RECT 83.650 120.250 83.970 120.310 ;
        RECT 93.785 120.265 94.075 120.310 ;
        RECT 97.925 120.265 98.215 120.310 ;
        RECT 105.270 120.250 105.590 120.310 ;
        RECT 106.205 120.450 106.495 120.495 ;
        RECT 109.195 120.450 109.730 120.495 ;
        RECT 106.205 120.310 109.730 120.450 ;
        RECT 106.205 120.265 106.495 120.310 ;
        RECT 109.195 120.265 109.730 120.310 ;
        RECT 109.410 120.250 109.730 120.265 ;
        RECT 109.960 120.310 118.840 120.450 ;
        RECT 34.400 120.110 34.690 120.155 ;
        RECT 34.400 119.970 36.935 120.110 ;
        RECT 34.400 119.925 34.690 119.970 ;
        RECT 22.025 119.770 22.315 119.815 ;
        RECT 30.750 119.770 31.070 119.830 ;
        RECT 22.025 119.630 31.070 119.770 ;
        RECT 22.025 119.585 22.315 119.630 ;
        RECT 30.750 119.570 31.070 119.630 ;
        RECT 32.540 119.770 32.830 119.815 ;
        RECT 34.890 119.770 35.210 119.830 ;
        RECT 36.720 119.815 36.935 119.970 ;
        RECT 37.650 119.910 37.970 120.170 ;
        RECT 39.505 119.925 39.795 120.155 ;
        RECT 35.800 119.770 36.090 119.815 ;
        RECT 32.540 119.630 36.090 119.770 ;
        RECT 32.540 119.585 32.830 119.630 ;
        RECT 34.890 119.570 35.210 119.630 ;
        RECT 35.800 119.585 36.090 119.630 ;
        RECT 36.720 119.770 37.010 119.815 ;
        RECT 38.580 119.770 38.870 119.815 ;
        RECT 36.720 119.630 38.870 119.770 ;
        RECT 39.580 119.770 39.720 119.925 ;
        RECT 41.790 119.910 42.110 120.170 ;
        RECT 45.470 119.910 45.790 120.170 ;
        RECT 46.480 120.110 46.620 120.250 ;
        RECT 47.785 120.110 48.075 120.155 ;
        RECT 46.480 119.970 48.075 120.110 ;
        RECT 47.785 119.925 48.075 119.970 ;
        RECT 50.070 120.110 50.390 120.170 ;
        RECT 50.545 120.110 50.835 120.155 ;
        RECT 54.225 120.110 54.515 120.155 ;
        RECT 50.070 119.970 54.515 120.110 ;
        RECT 50.070 119.910 50.390 119.970 ;
        RECT 50.545 119.925 50.835 119.970 ;
        RECT 54.225 119.925 54.515 119.970 ;
        RECT 55.605 120.110 55.895 120.155 ;
        RECT 57.890 120.110 58.210 120.170 ;
        RECT 55.605 119.970 58.210 120.110 ;
        RECT 55.605 119.925 55.895 119.970 ;
        RECT 57.890 119.910 58.210 119.970 ;
        RECT 63.380 120.110 63.670 120.155 ;
        RECT 63.380 119.970 65.915 120.110 ;
        RECT 63.380 119.925 63.670 119.970 ;
        RECT 46.390 119.770 46.710 119.830 ;
        RECT 39.580 119.630 46.710 119.770 ;
        RECT 36.720 119.585 37.010 119.630 ;
        RECT 38.580 119.585 38.870 119.630 ;
        RECT 46.390 119.570 46.710 119.630 ;
        RECT 61.520 119.770 61.810 119.815 ;
        RECT 62.030 119.770 62.350 119.830 ;
        RECT 65.700 119.815 65.915 119.970 ;
        RECT 68.485 119.925 68.775 120.155 ;
        RECT 64.780 119.770 65.070 119.815 ;
        RECT 61.520 119.630 65.070 119.770 ;
        RECT 61.520 119.585 61.810 119.630 ;
        RECT 62.030 119.570 62.350 119.630 ;
        RECT 64.780 119.585 65.070 119.630 ;
        RECT 65.700 119.770 65.990 119.815 ;
        RECT 67.560 119.770 67.850 119.815 ;
        RECT 65.700 119.630 67.850 119.770 ;
        RECT 68.560 119.770 68.700 119.925 ;
        RECT 69.850 119.910 70.170 120.170 ;
        RECT 73.070 120.110 73.390 120.170 ;
        RECT 74.465 120.110 74.755 120.155 ;
        RECT 81.825 120.110 82.115 120.155 ;
        RECT 73.070 119.970 74.755 120.110 ;
        RECT 73.070 119.910 73.390 119.970 ;
        RECT 74.465 119.925 74.755 119.970 ;
        RECT 80.520 119.970 82.115 120.110 ;
        RECT 70.770 119.770 71.090 119.830 ;
        RECT 68.560 119.630 71.090 119.770 ;
        RECT 65.700 119.585 65.990 119.630 ;
        RECT 67.560 119.585 67.850 119.630 ;
        RECT 70.770 119.570 71.090 119.630 ;
        RECT 78.145 119.770 78.435 119.815 ;
        RECT 79.510 119.770 79.830 119.830 ;
        RECT 78.145 119.630 79.830 119.770 ;
        RECT 78.145 119.585 78.435 119.630 ;
        RECT 79.510 119.570 79.830 119.630 ;
        RECT 20.185 119.430 20.475 119.475 ;
        RECT 21.090 119.430 21.410 119.490 ;
        RECT 20.185 119.290 21.410 119.430 ;
        RECT 20.185 119.245 20.475 119.290 ;
        RECT 21.090 119.230 21.410 119.290 ;
        RECT 25.230 119.430 25.550 119.490 ;
        RECT 26.165 119.430 26.455 119.475 ;
        RECT 25.230 119.290 26.455 119.430 ;
        RECT 25.230 119.230 25.550 119.290 ;
        RECT 26.165 119.245 26.455 119.290 ;
        RECT 39.950 119.230 40.270 119.490 ;
        RECT 42.250 119.230 42.570 119.490 ;
        RECT 44.565 119.430 44.855 119.475 ;
        RECT 45.010 119.430 45.330 119.490 ;
        RECT 44.565 119.290 45.330 119.430 ;
        RECT 44.565 119.245 44.855 119.290 ;
        RECT 45.010 119.230 45.330 119.290 ;
        RECT 49.610 119.230 49.930 119.490 ;
        RECT 50.990 119.230 51.310 119.490 ;
        RECT 74.925 119.430 75.215 119.475 ;
        RECT 75.370 119.430 75.690 119.490 ;
        RECT 74.925 119.290 75.690 119.430 ;
        RECT 74.925 119.245 75.215 119.290 ;
        RECT 75.370 119.230 75.690 119.290 ;
        RECT 78.605 119.430 78.895 119.475 ;
        RECT 79.050 119.430 79.370 119.490 ;
        RECT 80.520 119.475 80.660 119.970 ;
        RECT 81.825 119.925 82.115 119.970 ;
        RECT 83.190 119.910 83.510 120.170 ;
        RECT 84.110 119.910 84.430 120.170 ;
        RECT 93.310 120.110 93.630 120.170 ;
        RECT 99.290 120.110 99.610 120.170 ;
        RECT 93.310 119.970 99.610 120.110 ;
        RECT 93.310 119.910 93.630 119.970 ;
        RECT 99.290 119.910 99.610 119.970 ;
        RECT 100.210 120.110 100.530 120.170 ;
        RECT 103.445 120.110 103.735 120.155 ;
        RECT 109.960 120.110 110.100 120.310 ;
        RECT 118.700 120.170 118.840 120.310 ;
        RECT 100.210 119.970 110.100 120.110 ;
        RECT 113.060 120.110 113.350 120.155 ;
        RECT 113.060 119.970 115.595 120.110 ;
        RECT 100.210 119.910 100.530 119.970 ;
        RECT 103.445 119.925 103.735 119.970 ;
        RECT 113.060 119.925 113.350 119.970 ;
        RECT 98.845 119.770 99.135 119.815 ;
        RECT 102.510 119.770 102.830 119.830 ;
        RECT 106.190 119.770 106.510 119.830 ;
        RECT 106.665 119.770 106.955 119.815 ;
        RECT 98.845 119.630 106.955 119.770 ;
        RECT 98.845 119.585 99.135 119.630 ;
        RECT 102.510 119.570 102.830 119.630 ;
        RECT 106.190 119.570 106.510 119.630 ;
        RECT 106.665 119.585 106.955 119.630 ;
        RECT 111.200 119.770 111.490 119.815 ;
        RECT 113.550 119.770 113.870 119.830 ;
        RECT 115.380 119.815 115.595 119.970 ;
        RECT 116.310 119.910 116.630 120.170 ;
        RECT 118.165 119.925 118.455 120.155 ;
        RECT 114.460 119.770 114.750 119.815 ;
        RECT 111.200 119.630 114.750 119.770 ;
        RECT 111.200 119.585 111.490 119.630 ;
        RECT 113.550 119.570 113.870 119.630 ;
        RECT 114.460 119.585 114.750 119.630 ;
        RECT 115.380 119.770 115.670 119.815 ;
        RECT 117.240 119.770 117.530 119.815 ;
        RECT 115.380 119.630 117.530 119.770 ;
        RECT 115.380 119.585 115.670 119.630 ;
        RECT 117.240 119.585 117.530 119.630 ;
        RECT 78.605 119.290 79.370 119.430 ;
        RECT 78.605 119.245 78.895 119.290 ;
        RECT 79.050 119.230 79.370 119.290 ;
        RECT 80.445 119.245 80.735 119.475 ;
        RECT 80.890 119.230 81.210 119.490 ;
        RECT 82.730 119.230 83.050 119.490 ;
        RECT 84.570 119.430 84.890 119.490 ;
        RECT 85.045 119.430 85.335 119.475 ;
        RECT 84.570 119.290 85.335 119.430 ;
        RECT 84.570 119.230 84.890 119.290 ;
        RECT 85.045 119.245 85.335 119.290 ;
        RECT 87.330 119.430 87.650 119.490 ;
        RECT 91.025 119.430 91.315 119.475 ;
        RECT 87.330 119.290 91.315 119.430 ;
        RECT 87.330 119.230 87.650 119.290 ;
        RECT 91.025 119.245 91.315 119.290 ;
        RECT 92.865 119.430 93.155 119.475 ;
        RECT 93.770 119.430 94.090 119.490 ;
        RECT 92.865 119.290 94.090 119.430 ;
        RECT 92.865 119.245 93.155 119.290 ;
        RECT 93.770 119.230 94.090 119.290 ;
        RECT 101.130 119.230 101.450 119.490 ;
        RECT 103.905 119.430 104.195 119.475 ;
        RECT 105.730 119.430 106.050 119.490 ;
        RECT 103.905 119.290 106.050 119.430 ;
        RECT 103.905 119.245 104.195 119.290 ;
        RECT 105.730 119.230 106.050 119.290 ;
        RECT 108.505 119.430 108.795 119.475 ;
        RECT 108.950 119.430 109.270 119.490 ;
        RECT 108.505 119.290 109.270 119.430 ;
        RECT 108.505 119.245 108.795 119.290 ;
        RECT 108.950 119.230 109.270 119.290 ;
        RECT 111.710 119.430 112.030 119.490 ;
        RECT 118.240 119.430 118.380 119.925 ;
        RECT 118.610 119.910 118.930 120.170 ;
        RECT 120.450 119.910 120.770 120.170 ;
        RECT 111.710 119.290 118.380 119.430 ;
        RECT 111.710 119.230 112.030 119.290 ;
        RECT 14.580 118.610 127.740 119.090 ;
        RECT 18.115 118.410 18.405 118.455 ;
        RECT 22.470 118.410 22.790 118.470 ;
        RECT 18.115 118.270 22.790 118.410 ;
        RECT 18.115 118.225 18.405 118.270 ;
        RECT 22.470 118.210 22.790 118.270 ;
        RECT 36.270 118.455 36.590 118.470 ;
        RECT 36.270 118.225 36.805 118.455 ;
        RECT 37.895 118.410 38.185 118.455 ;
        RECT 42.250 118.410 42.570 118.470 ;
        RECT 37.895 118.270 42.570 118.410 ;
        RECT 37.895 118.225 38.185 118.270 ;
        RECT 36.270 118.210 36.590 118.225 ;
        RECT 42.250 118.210 42.570 118.270 ;
        RECT 62.030 118.210 62.350 118.470 ;
        RECT 63.655 118.410 63.945 118.455 ;
        RECT 64.330 118.410 64.650 118.470 ;
        RECT 63.655 118.270 64.650 118.410 ;
        RECT 63.655 118.225 63.945 118.270 ;
        RECT 64.330 118.210 64.650 118.270 ;
        RECT 73.315 118.410 73.605 118.455 ;
        RECT 79.050 118.410 79.370 118.470 ;
        RECT 73.315 118.270 79.370 118.410 ;
        RECT 73.315 118.225 73.605 118.270 ;
        RECT 79.050 118.210 79.370 118.270 ;
        RECT 82.745 118.410 83.035 118.455 ;
        RECT 84.110 118.410 84.430 118.470 ;
        RECT 93.310 118.455 93.630 118.470 ;
        RECT 82.745 118.270 84.430 118.410 ;
        RECT 82.745 118.225 83.035 118.270 ;
        RECT 84.110 118.210 84.430 118.270 ;
        RECT 93.095 118.225 93.630 118.455 ;
        RECT 93.310 118.210 93.630 118.225 ;
        RECT 102.510 118.455 102.830 118.470 ;
        RECT 102.510 118.225 103.045 118.455 ;
        RECT 102.510 118.210 102.830 118.225 ;
        RECT 113.550 118.210 113.870 118.470 ;
        RECT 116.310 118.210 116.630 118.470 ;
        RECT 23.390 118.115 23.710 118.130 ;
        RECT 20.120 118.070 20.410 118.115 ;
        RECT 23.380 118.070 23.710 118.115 ;
        RECT 20.120 117.930 23.710 118.070 ;
        RECT 20.120 117.885 20.410 117.930 ;
        RECT 23.380 117.885 23.710 117.930 ;
        RECT 23.390 117.870 23.710 117.885 ;
        RECT 24.300 118.070 24.590 118.115 ;
        RECT 26.160 118.070 26.450 118.115 ;
        RECT 24.300 117.930 26.450 118.070 ;
        RECT 24.300 117.885 24.590 117.930 ;
        RECT 26.160 117.885 26.450 117.930 ;
        RECT 28.470 118.070 28.760 118.115 ;
        RECT 30.330 118.070 30.620 118.115 ;
        RECT 28.470 117.930 30.620 118.070 ;
        RECT 28.470 117.885 28.760 117.930 ;
        RECT 30.330 117.885 30.620 117.930 ;
        RECT 31.250 118.070 31.540 118.115 ;
        RECT 34.510 118.070 34.800 118.115 ;
        RECT 35.350 118.070 35.670 118.130 ;
        RECT 43.170 118.115 43.490 118.130 ;
        RECT 31.250 117.930 35.670 118.070 ;
        RECT 31.250 117.885 31.540 117.930 ;
        RECT 34.510 117.885 34.800 117.930 ;
        RECT 17.425 117.730 17.715 117.775 ;
        RECT 19.250 117.730 19.570 117.790 ;
        RECT 17.425 117.590 19.570 117.730 ;
        RECT 17.425 117.545 17.715 117.590 ;
        RECT 19.250 117.530 19.570 117.590 ;
        RECT 21.980 117.730 22.270 117.775 ;
        RECT 24.300 117.730 24.515 117.885 ;
        RECT 21.980 117.590 24.515 117.730 ;
        RECT 21.980 117.545 22.270 117.590 ;
        RECT 25.230 117.530 25.550 117.790 ;
        RECT 30.405 117.730 30.620 117.885 ;
        RECT 35.350 117.870 35.670 117.930 ;
        RECT 39.900 118.070 40.190 118.115 ;
        RECT 43.160 118.070 43.490 118.115 ;
        RECT 39.900 117.930 43.490 118.070 ;
        RECT 39.900 117.885 40.190 117.930 ;
        RECT 43.160 117.885 43.490 117.930 ;
        RECT 43.170 117.870 43.490 117.885 ;
        RECT 44.080 118.070 44.370 118.115 ;
        RECT 45.940 118.070 46.230 118.115 ;
        RECT 44.080 117.930 46.230 118.070 ;
        RECT 44.080 117.885 44.370 117.930 ;
        RECT 45.940 117.885 46.230 117.930 ;
        RECT 49.560 118.070 49.850 118.115 ;
        RECT 50.990 118.070 51.310 118.130 ;
        RECT 52.820 118.070 53.110 118.115 ;
        RECT 49.560 117.930 53.110 118.070 ;
        RECT 49.560 117.885 49.850 117.930 ;
        RECT 32.650 117.730 32.940 117.775 ;
        RECT 30.405 117.590 32.940 117.730 ;
        RECT 32.650 117.545 32.940 117.590 ;
        RECT 41.760 117.730 42.050 117.775 ;
        RECT 44.080 117.730 44.295 117.885 ;
        RECT 50.990 117.870 51.310 117.930 ;
        RECT 52.820 117.885 53.110 117.930 ;
        RECT 53.740 118.070 54.030 118.115 ;
        RECT 55.600 118.070 55.890 118.115 ;
        RECT 53.740 117.930 55.890 118.070 ;
        RECT 53.740 117.885 54.030 117.930 ;
        RECT 55.600 117.885 55.890 117.930 ;
        RECT 65.660 118.070 65.950 118.115 ;
        RECT 66.630 118.070 66.950 118.130 ;
        RECT 75.370 118.115 75.690 118.130 ;
        RECT 68.920 118.070 69.210 118.115 ;
        RECT 65.660 117.930 69.210 118.070 ;
        RECT 65.660 117.885 65.950 117.930 ;
        RECT 41.760 117.590 44.295 117.730 ;
        RECT 41.760 117.545 42.050 117.590 ;
        RECT 45.010 117.530 45.330 117.790 ;
        RECT 46.390 117.730 46.710 117.790 ;
        RECT 46.865 117.730 47.155 117.775 ;
        RECT 46.390 117.590 47.155 117.730 ;
        RECT 46.390 117.530 46.710 117.590 ;
        RECT 46.865 117.545 47.155 117.590 ;
        RECT 51.420 117.730 51.710 117.775 ;
        RECT 53.740 117.730 53.955 117.885 ;
        RECT 66.630 117.870 66.950 117.930 ;
        RECT 68.920 117.885 69.210 117.930 ;
        RECT 69.840 118.070 70.130 118.115 ;
        RECT 71.700 118.070 71.990 118.115 ;
        RECT 69.840 117.930 71.990 118.070 ;
        RECT 69.840 117.885 70.130 117.930 ;
        RECT 71.700 117.885 71.990 117.930 ;
        RECT 75.320 118.070 75.690 118.115 ;
        RECT 78.580 118.070 78.870 118.115 ;
        RECT 75.320 117.930 78.870 118.070 ;
        RECT 75.320 117.885 75.690 117.930 ;
        RECT 78.580 117.885 78.870 117.930 ;
        RECT 79.500 118.070 79.790 118.115 ;
        RECT 81.360 118.070 81.650 118.115 ;
        RECT 79.500 117.930 81.650 118.070 ;
        RECT 79.500 117.885 79.790 117.930 ;
        RECT 81.360 117.885 81.650 117.930 ;
        RECT 83.190 118.070 83.510 118.130 ;
        RECT 89.645 118.070 89.935 118.115 ;
        RECT 95.100 118.070 95.390 118.115 ;
        RECT 98.360 118.070 98.650 118.115 ;
        RECT 83.190 117.930 89.400 118.070 ;
        RECT 51.420 117.590 53.955 117.730 ;
        RECT 51.420 117.545 51.710 117.590 ;
        RECT 25.690 117.390 26.010 117.450 ;
        RECT 27.085 117.390 27.375 117.435 ;
        RECT 27.545 117.390 27.835 117.435 ;
        RECT 25.690 117.250 27.835 117.390 ;
        RECT 25.690 117.190 26.010 117.250 ;
        RECT 27.085 117.205 27.375 117.250 ;
        RECT 27.545 117.205 27.835 117.250 ;
        RECT 29.385 117.390 29.675 117.435 ;
        RECT 39.030 117.390 39.350 117.450 ;
        RECT 29.385 117.250 39.350 117.390 ;
        RECT 46.940 117.390 47.080 117.545 ;
        RECT 54.670 117.530 54.990 117.790 ;
        RECT 57.890 117.730 58.210 117.790 ;
        RECT 59.730 117.730 60.050 117.790 ;
        RECT 61.585 117.730 61.875 117.775 ;
        RECT 57.890 117.590 61.875 117.730 ;
        RECT 57.890 117.530 58.210 117.590 ;
        RECT 59.730 117.530 60.050 117.590 ;
        RECT 61.585 117.545 61.875 117.590 ;
        RECT 67.520 117.730 67.810 117.775 ;
        RECT 69.840 117.730 70.055 117.885 ;
        RECT 75.370 117.870 75.690 117.885 ;
        RECT 67.520 117.590 70.055 117.730 ;
        RECT 77.180 117.730 77.470 117.775 ;
        RECT 79.500 117.730 79.715 117.885 ;
        RECT 83.190 117.870 83.510 117.930 ;
        RECT 77.180 117.590 79.715 117.730 ;
        RECT 80.445 117.730 80.735 117.775 ;
        RECT 80.890 117.730 81.210 117.790 ;
        RECT 84.585 117.730 84.875 117.775 ;
        RECT 80.445 117.590 81.210 117.730 ;
        RECT 67.520 117.545 67.810 117.590 ;
        RECT 77.180 117.545 77.470 117.590 ;
        RECT 80.445 117.545 80.735 117.590 ;
        RECT 56.510 117.390 56.830 117.450 ;
        RECT 46.940 117.250 56.830 117.390 ;
        RECT 61.660 117.390 61.800 117.545 ;
        RECT 80.890 117.530 81.210 117.590 ;
        RECT 81.440 117.590 84.875 117.730 ;
        RECT 69.390 117.390 69.710 117.450 ;
        RECT 61.660 117.250 69.710 117.390 ;
        RECT 29.385 117.205 29.675 117.250 ;
        RECT 39.030 117.190 39.350 117.250 ;
        RECT 56.510 117.190 56.830 117.250 ;
        RECT 69.390 117.190 69.710 117.250 ;
        RECT 70.770 117.190 71.090 117.450 ;
        RECT 71.230 117.390 71.550 117.450 ;
        RECT 72.625 117.390 72.915 117.435 ;
        RECT 71.230 117.250 72.915 117.390 ;
        RECT 71.230 117.190 71.550 117.250 ;
        RECT 72.625 117.205 72.915 117.250 ;
        RECT 79.510 117.390 79.830 117.450 ;
        RECT 81.440 117.390 81.580 117.590 ;
        RECT 84.585 117.545 84.875 117.590 ;
        RECT 85.045 117.730 85.335 117.775 ;
        RECT 85.045 117.590 87.100 117.730 ;
        RECT 85.045 117.545 85.335 117.590 ;
        RECT 79.510 117.250 81.580 117.390 ;
        RECT 82.285 117.390 82.575 117.435 ;
        RECT 85.490 117.390 85.810 117.450 ;
        RECT 82.285 117.250 85.810 117.390 ;
        RECT 79.510 117.190 79.830 117.250 ;
        RECT 82.285 117.205 82.575 117.250 ;
        RECT 85.490 117.190 85.810 117.250 ;
        RECT 85.965 117.205 86.255 117.435 ;
        RECT 86.960 117.390 87.100 117.590 ;
        RECT 87.330 117.530 87.650 117.790 ;
        RECT 89.260 117.775 89.400 117.930 ;
        RECT 89.645 117.930 98.650 118.070 ;
        RECT 89.645 117.885 89.935 117.930 ;
        RECT 95.100 117.885 95.390 117.930 ;
        RECT 98.360 117.885 98.650 117.930 ;
        RECT 99.280 118.070 99.570 118.115 ;
        RECT 101.140 118.070 101.430 118.115 ;
        RECT 99.280 117.930 101.430 118.070 ;
        RECT 99.280 117.885 99.570 117.930 ;
        RECT 101.140 117.885 101.430 117.930 ;
        RECT 104.760 118.070 105.050 118.115 ;
        RECT 105.730 118.070 106.050 118.130 ;
        RECT 108.020 118.070 108.310 118.115 ;
        RECT 104.760 117.930 108.310 118.070 ;
        RECT 104.760 117.885 105.050 117.930 ;
        RECT 89.185 117.730 89.475 117.775 ;
        RECT 90.565 117.730 90.855 117.775 ;
        RECT 89.185 117.590 90.855 117.730 ;
        RECT 89.185 117.545 89.475 117.590 ;
        RECT 90.565 117.545 90.855 117.590 ;
        RECT 96.960 117.730 97.250 117.775 ;
        RECT 99.280 117.730 99.495 117.885 ;
        RECT 105.730 117.870 106.050 117.930 ;
        RECT 108.020 117.885 108.310 117.930 ;
        RECT 108.940 118.070 109.230 118.115 ;
        RECT 110.800 118.070 111.090 118.115 ;
        RECT 118.150 118.070 118.470 118.130 ;
        RECT 108.940 117.930 111.090 118.070 ;
        RECT 108.940 117.885 109.230 117.930 ;
        RECT 110.800 117.885 111.090 117.930 ;
        RECT 114.100 117.930 118.470 118.070 ;
        RECT 96.960 117.590 99.495 117.730 ;
        RECT 106.620 117.730 106.910 117.775 ;
        RECT 108.940 117.730 109.155 117.885 ;
        RECT 106.620 117.590 109.155 117.730 ;
        RECT 96.960 117.545 97.250 117.590 ;
        RECT 106.620 117.545 106.910 117.590 ;
        RECT 109.870 117.530 110.190 117.790 ;
        RECT 111.710 117.530 112.030 117.790 ;
        RECT 114.100 117.775 114.240 117.930 ;
        RECT 118.150 117.870 118.470 117.930 ;
        RECT 114.025 117.545 114.315 117.775 ;
        RECT 115.390 117.530 115.710 117.790 ;
        RECT 93.770 117.390 94.090 117.450 ;
        RECT 86.960 117.250 94.090 117.390 ;
        RECT 21.980 117.050 22.270 117.095 ;
        RECT 24.760 117.050 25.050 117.095 ;
        RECT 26.620 117.050 26.910 117.095 ;
        RECT 21.980 116.910 26.910 117.050 ;
        RECT 21.980 116.865 22.270 116.910 ;
        RECT 24.760 116.865 25.050 116.910 ;
        RECT 26.620 116.865 26.910 116.910 ;
        RECT 28.010 117.050 28.300 117.095 ;
        RECT 29.870 117.050 30.160 117.095 ;
        RECT 32.650 117.050 32.940 117.095 ;
        RECT 28.010 116.910 32.940 117.050 ;
        RECT 28.010 116.865 28.300 116.910 ;
        RECT 29.870 116.865 30.160 116.910 ;
        RECT 32.650 116.865 32.940 116.910 ;
        RECT 41.760 117.050 42.050 117.095 ;
        RECT 44.540 117.050 44.830 117.095 ;
        RECT 46.400 117.050 46.690 117.095 ;
        RECT 41.760 116.910 46.690 117.050 ;
        RECT 41.760 116.865 42.050 116.910 ;
        RECT 44.540 116.865 44.830 116.910 ;
        RECT 46.400 116.865 46.690 116.910 ;
        RECT 51.420 117.050 51.710 117.095 ;
        RECT 54.200 117.050 54.490 117.095 ;
        RECT 56.060 117.050 56.350 117.095 ;
        RECT 51.420 116.910 56.350 117.050 ;
        RECT 51.420 116.865 51.710 116.910 ;
        RECT 54.200 116.865 54.490 116.910 ;
        RECT 56.060 116.865 56.350 116.910 ;
        RECT 67.520 117.050 67.810 117.095 ;
        RECT 70.300 117.050 70.590 117.095 ;
        RECT 72.160 117.050 72.450 117.095 ;
        RECT 67.520 116.910 72.450 117.050 ;
        RECT 67.520 116.865 67.810 116.910 ;
        RECT 70.300 116.865 70.590 116.910 ;
        RECT 72.160 116.865 72.450 116.910 ;
        RECT 77.180 117.050 77.470 117.095 ;
        RECT 79.960 117.050 80.250 117.095 ;
        RECT 81.820 117.050 82.110 117.095 ;
        RECT 77.180 116.910 82.110 117.050 ;
        RECT 77.180 116.865 77.470 116.910 ;
        RECT 79.960 116.865 80.250 116.910 ;
        RECT 81.820 116.865 82.110 116.910 ;
        RECT 83.650 117.050 83.970 117.110 ;
        RECT 86.040 117.050 86.180 117.205 ;
        RECT 93.770 117.190 94.090 117.250 ;
        RECT 100.210 117.190 100.530 117.450 ;
        RECT 102.065 117.390 102.355 117.435 ;
        RECT 111.800 117.390 111.940 117.530 ;
        RECT 102.065 117.250 111.940 117.390 ;
        RECT 102.065 117.205 102.355 117.250 ;
        RECT 83.650 116.910 86.180 117.050 ;
        RECT 96.960 117.050 97.250 117.095 ;
        RECT 99.740 117.050 100.030 117.095 ;
        RECT 101.600 117.050 101.890 117.095 ;
        RECT 96.960 116.910 101.890 117.050 ;
        RECT 83.650 116.850 83.970 116.910 ;
        RECT 96.960 116.865 97.250 116.910 ;
        RECT 99.740 116.865 100.030 116.910 ;
        RECT 101.600 116.865 101.890 116.910 ;
        RECT 106.620 117.050 106.910 117.095 ;
        RECT 109.400 117.050 109.690 117.095 ;
        RECT 111.260 117.050 111.550 117.095 ;
        RECT 106.620 116.910 111.550 117.050 ;
        RECT 106.620 116.865 106.910 116.910 ;
        RECT 109.400 116.865 109.690 116.910 ;
        RECT 111.260 116.865 111.550 116.910 ;
        RECT 16.965 116.710 17.255 116.755 ;
        RECT 28.450 116.710 28.770 116.770 ;
        RECT 16.965 116.570 28.770 116.710 ;
        RECT 16.965 116.525 17.255 116.570 ;
        RECT 28.450 116.510 28.770 116.570 ;
        RECT 45.930 116.710 46.250 116.770 ;
        RECT 47.555 116.710 47.845 116.755 ;
        RECT 45.930 116.570 47.845 116.710 ;
        RECT 45.930 116.510 46.250 116.570 ;
        RECT 47.555 116.525 47.845 116.570 ;
        RECT 88.250 116.510 88.570 116.770 ;
        RECT 91.010 116.510 91.330 116.770 ;
        RECT 14.580 115.890 127.740 116.370 ;
        RECT 22.945 115.690 23.235 115.735 ;
        RECT 23.390 115.690 23.710 115.750 ;
        RECT 22.945 115.550 23.710 115.690 ;
        RECT 22.945 115.505 23.235 115.550 ;
        RECT 23.390 115.490 23.710 115.550 ;
        RECT 30.750 115.690 31.070 115.750 ;
        RECT 33.755 115.690 34.045 115.735 ;
        RECT 30.750 115.550 34.045 115.690 ;
        RECT 30.750 115.490 31.070 115.550 ;
        RECT 33.755 115.505 34.045 115.550 ;
        RECT 35.350 115.490 35.670 115.750 ;
        RECT 37.650 115.490 37.970 115.750 ;
        RECT 39.030 115.490 39.350 115.750 ;
        RECT 43.170 115.690 43.490 115.750 ;
        RECT 44.565 115.690 44.855 115.735 ;
        RECT 43.170 115.550 44.855 115.690 ;
        RECT 43.170 115.490 43.490 115.550 ;
        RECT 44.565 115.505 44.855 115.550 ;
        RECT 45.470 115.490 45.790 115.750 ;
        RECT 53.305 115.690 53.595 115.735 ;
        RECT 54.670 115.690 54.990 115.750 ;
        RECT 53.305 115.550 54.990 115.690 ;
        RECT 53.305 115.505 53.595 115.550 ;
        RECT 54.670 115.490 54.990 115.550 ;
        RECT 66.630 115.490 66.950 115.750 ;
        RECT 68.945 115.690 69.235 115.735 ;
        RECT 70.770 115.690 71.090 115.750 ;
        RECT 68.945 115.550 71.090 115.690 ;
        RECT 68.945 115.505 69.235 115.550 ;
        RECT 70.770 115.490 71.090 115.550 ;
        RECT 71.230 115.690 71.550 115.750 ;
        RECT 73.530 115.690 73.850 115.750 ;
        RECT 71.230 115.550 73.850 115.690 ;
        RECT 71.230 115.490 71.550 115.550 ;
        RECT 73.530 115.490 73.850 115.550 ;
        RECT 77.455 115.690 77.745 115.735 ;
        RECT 79.510 115.690 79.830 115.750 ;
        RECT 77.455 115.550 79.830 115.690 ;
        RECT 77.455 115.505 77.745 115.550 ;
        RECT 79.510 115.490 79.830 115.550 ;
        RECT 93.770 115.690 94.090 115.750 ;
        RECT 96.315 115.690 96.605 115.735 ;
        RECT 93.770 115.550 96.605 115.690 ;
        RECT 93.770 115.490 94.090 115.550 ;
        RECT 96.315 115.505 96.605 115.550 ;
        RECT 100.210 115.490 100.530 115.750 ;
        RECT 108.965 115.690 109.255 115.735 ;
        RECT 109.870 115.690 110.190 115.750 ;
        RECT 108.965 115.550 110.190 115.690 ;
        RECT 108.965 115.505 109.255 115.550 ;
        RECT 109.870 115.490 110.190 115.550 ;
        RECT 114.945 115.690 115.235 115.735 ;
        RECT 115.390 115.690 115.710 115.750 ;
        RECT 114.945 115.550 115.710 115.690 ;
        RECT 114.945 115.505 115.235 115.550 ;
        RECT 115.390 115.490 115.710 115.550 ;
        RECT 22.025 115.165 22.315 115.395 ;
        RECT 25.250 115.350 25.540 115.395 ;
        RECT 27.110 115.350 27.400 115.395 ;
        RECT 29.890 115.350 30.180 115.395 ;
        RECT 25.250 115.210 30.180 115.350 ;
        RECT 25.250 115.165 25.540 115.210 ;
        RECT 27.110 115.165 27.400 115.210 ;
        RECT 29.890 115.165 30.180 115.210 ;
        RECT 43.630 115.350 43.950 115.410 ;
        RECT 81.320 115.350 81.610 115.395 ;
        RECT 84.100 115.350 84.390 115.395 ;
        RECT 85.960 115.350 86.250 115.395 ;
        RECT 43.630 115.210 48.460 115.350 ;
        RECT 19.710 115.010 20.030 115.070 ;
        RECT 22.100 115.010 22.240 115.165 ;
        RECT 43.630 115.150 43.950 115.210 ;
        RECT 24.785 115.010 25.075 115.055 ;
        RECT 25.690 115.010 26.010 115.070 ;
        RECT 45.930 115.010 46.250 115.070 ;
        RECT 48.320 115.055 48.460 115.210 ;
        RECT 81.320 115.210 86.250 115.350 ;
        RECT 81.320 115.165 81.610 115.210 ;
        RECT 84.100 115.165 84.390 115.210 ;
        RECT 85.960 115.165 86.250 115.210 ;
        RECT 87.810 115.350 88.100 115.395 ;
        RECT 89.670 115.350 89.960 115.395 ;
        RECT 92.450 115.350 92.740 115.395 ;
        RECT 113.090 115.350 113.410 115.410 ;
        RECT 87.810 115.210 92.740 115.350 ;
        RECT 87.810 115.165 88.100 115.210 ;
        RECT 89.670 115.165 89.960 115.210 ;
        RECT 92.450 115.165 92.740 115.210 ;
        RECT 112.260 115.210 113.410 115.350 ;
        RECT 47.785 115.010 48.075 115.055 ;
        RECT 19.710 114.870 21.780 115.010 ;
        RECT 22.100 114.870 24.540 115.010 ;
        RECT 19.710 114.810 20.030 114.870 ;
        RECT 21.090 114.470 21.410 114.730 ;
        RECT 21.640 114.670 21.780 114.870 ;
        RECT 23.405 114.670 23.695 114.715 ;
        RECT 24.400 114.670 24.540 114.870 ;
        RECT 24.785 114.870 26.010 115.010 ;
        RECT 24.785 114.825 25.075 114.870 ;
        RECT 25.690 114.810 26.010 114.870 ;
        RECT 35.900 114.870 45.240 115.010 ;
        RECT 35.900 114.730 36.040 114.870 ;
        RECT 26.625 114.670 26.915 114.715 ;
        RECT 29.890 114.670 30.180 114.715 ;
        RECT 21.640 114.530 24.080 114.670 ;
        RECT 24.400 114.530 26.915 114.670 ;
        RECT 23.405 114.485 23.695 114.530 ;
        RECT 23.940 113.990 24.080 114.530 ;
        RECT 26.625 114.485 26.915 114.530 ;
        RECT 27.645 114.530 30.180 114.670 ;
        RECT 27.645 114.375 27.860 114.530 ;
        RECT 29.890 114.485 30.180 114.530 ;
        RECT 35.810 114.470 36.130 114.730 ;
        RECT 36.730 114.470 37.050 114.730 ;
        RECT 39.950 114.470 40.270 114.730 ;
        RECT 45.100 114.715 45.240 114.870 ;
        RECT 45.930 114.870 48.075 115.010 ;
        RECT 45.930 114.810 46.250 114.870 ;
        RECT 47.785 114.825 48.075 114.870 ;
        RECT 48.245 114.825 48.535 115.055 ;
        RECT 50.070 115.010 50.390 115.070 ;
        RECT 69.390 115.010 69.710 115.070 ;
        RECT 49.240 114.870 50.390 115.010 ;
        RECT 45.025 114.670 45.315 114.715 ;
        RECT 49.240 114.670 49.380 114.870 ;
        RECT 50.070 114.810 50.390 114.870 ;
        RECT 66.260 114.870 69.710 115.010 ;
        RECT 45.025 114.530 49.380 114.670 ;
        RECT 49.610 114.670 49.930 114.730 ;
        RECT 66.260 114.715 66.400 114.870 ;
        RECT 69.390 114.810 69.710 114.870 ;
        RECT 84.570 114.810 84.890 115.070 ;
        RECT 85.490 115.010 85.810 115.070 ;
        RECT 86.410 115.010 86.730 115.070 ;
        RECT 87.345 115.010 87.635 115.055 ;
        RECT 85.490 114.870 87.635 115.010 ;
        RECT 85.490 114.810 85.810 114.870 ;
        RECT 86.410 114.810 86.730 114.870 ;
        RECT 87.345 114.825 87.635 114.870 ;
        RECT 88.250 115.010 88.570 115.070 ;
        RECT 112.260 115.055 112.400 115.210 ;
        RECT 113.090 115.150 113.410 115.210 ;
        RECT 89.185 115.010 89.475 115.055 ;
        RECT 88.250 114.870 89.475 115.010 ;
        RECT 88.250 114.810 88.570 114.870 ;
        RECT 89.185 114.825 89.475 114.870 ;
        RECT 112.185 114.825 112.475 115.055 ;
        RECT 112.630 114.810 112.950 115.070 ;
        RECT 52.385 114.670 52.675 114.715 ;
        RECT 49.610 114.530 52.675 114.670 ;
        RECT 45.025 114.485 45.315 114.530 ;
        RECT 49.610 114.470 49.930 114.530 ;
        RECT 52.385 114.485 52.675 114.530 ;
        RECT 66.185 114.485 66.475 114.715 ;
        RECT 68.010 114.470 68.330 114.730 ;
        RECT 81.320 114.670 81.610 114.715 ;
        RECT 92.450 114.670 92.740 114.715 ;
        RECT 81.320 114.530 83.855 114.670 ;
        RECT 81.320 114.485 81.610 114.530 ;
        RECT 25.710 114.330 26.000 114.375 ;
        RECT 27.570 114.330 27.860 114.375 ;
        RECT 25.710 114.190 27.860 114.330 ;
        RECT 25.710 114.145 26.000 114.190 ;
        RECT 27.570 114.145 27.860 114.190 ;
        RECT 28.450 114.375 28.770 114.390 ;
        RECT 28.450 114.330 28.780 114.375 ;
        RECT 31.750 114.330 32.040 114.375 ;
        RECT 28.450 114.190 32.040 114.330 ;
        RECT 28.450 114.145 28.780 114.190 ;
        RECT 31.750 114.145 32.040 114.190 ;
        RECT 42.250 114.330 42.570 114.390 ;
        RECT 82.730 114.375 83.050 114.390 ;
        RECT 47.325 114.330 47.615 114.375 ;
        RECT 42.250 114.190 47.615 114.330 ;
        RECT 28.450 114.130 28.770 114.145 ;
        RECT 42.250 114.130 42.570 114.190 ;
        RECT 47.325 114.145 47.615 114.190 ;
        RECT 79.460 114.330 79.750 114.375 ;
        RECT 82.720 114.330 83.050 114.375 ;
        RECT 79.460 114.190 83.050 114.330 ;
        RECT 79.460 114.145 79.750 114.190 ;
        RECT 82.720 114.145 83.050 114.190 ;
        RECT 83.640 114.375 83.855 114.530 ;
        RECT 90.205 114.530 92.740 114.670 ;
        RECT 90.205 114.375 90.420 114.530 ;
        RECT 92.450 114.485 92.740 114.530 ;
        RECT 101.130 114.470 101.450 114.730 ;
        RECT 108.045 114.670 108.335 114.715 ;
        RECT 108.950 114.670 109.270 114.730 ;
        RECT 108.045 114.530 109.270 114.670 ;
        RECT 108.045 114.485 108.335 114.530 ;
        RECT 108.950 114.470 109.270 114.530 ;
        RECT 109.410 114.670 109.730 114.730 ;
        RECT 113.105 114.670 113.395 114.715 ;
        RECT 109.410 114.530 113.395 114.670 ;
        RECT 109.410 114.470 109.730 114.530 ;
        RECT 113.105 114.485 113.395 114.530 ;
        RECT 83.640 114.330 83.930 114.375 ;
        RECT 85.500 114.330 85.790 114.375 ;
        RECT 83.640 114.190 85.790 114.330 ;
        RECT 83.640 114.145 83.930 114.190 ;
        RECT 85.500 114.145 85.790 114.190 ;
        RECT 88.270 114.330 88.560 114.375 ;
        RECT 90.130 114.330 90.420 114.375 ;
        RECT 88.270 114.190 90.420 114.330 ;
        RECT 88.270 114.145 88.560 114.190 ;
        RECT 90.130 114.145 90.420 114.190 ;
        RECT 91.010 114.375 91.330 114.390 ;
        RECT 91.010 114.330 91.340 114.375 ;
        RECT 94.310 114.330 94.600 114.375 ;
        RECT 91.010 114.190 94.600 114.330 ;
        RECT 91.010 114.145 91.340 114.190 ;
        RECT 94.310 114.145 94.600 114.190 ;
        RECT 82.730 114.130 83.050 114.145 ;
        RECT 91.010 114.130 91.330 114.145 ;
        RECT 35.810 113.990 36.130 114.050 ;
        RECT 23.940 113.850 36.130 113.990 ;
        RECT 35.810 113.790 36.130 113.850 ;
        RECT 101.590 113.990 101.910 114.050 ;
        RECT 121.830 113.990 122.150 114.050 ;
        RECT 101.590 113.850 122.150 113.990 ;
        RECT 101.590 113.790 101.910 113.850 ;
        RECT 121.830 113.790 122.150 113.850 ;
        RECT 14.580 113.170 127.740 113.650 ;
        RECT 34.445 112.970 34.735 113.015 ;
        RECT 34.890 112.970 35.210 113.030 ;
        RECT 34.445 112.830 35.210 112.970 ;
        RECT 34.445 112.785 34.735 112.830 ;
        RECT 34.890 112.770 35.210 112.830 ;
        RECT 102.985 112.970 103.275 113.015 ;
        RECT 111.710 112.970 112.030 113.030 ;
        RECT 102.985 112.830 112.030 112.970 ;
        RECT 102.985 112.785 103.275 112.830 ;
        RECT 18.905 112.630 19.195 112.675 ;
        RECT 21.090 112.630 21.410 112.690 ;
        RECT 22.145 112.630 22.795 112.675 ;
        RECT 18.905 112.490 22.795 112.630 ;
        RECT 18.905 112.445 19.495 112.490 ;
        RECT 19.205 112.130 19.495 112.445 ;
        RECT 21.090 112.430 21.410 112.490 ;
        RECT 22.145 112.445 22.795 112.490 ;
        RECT 46.865 112.630 47.155 112.675 ;
        RECT 49.150 112.630 49.470 112.690 ;
        RECT 46.865 112.490 49.470 112.630 ;
        RECT 46.865 112.445 47.155 112.490 ;
        RECT 49.150 112.430 49.470 112.490 ;
        RECT 92.850 112.430 93.170 112.690 ;
        RECT 101.605 112.630 101.895 112.675 ;
        RECT 103.060 112.630 103.200 112.785 ;
        RECT 111.710 112.770 112.030 112.830 ;
        RECT 117.230 112.970 117.550 113.030 ;
        RECT 120.925 112.970 121.215 113.015 ;
        RECT 117.230 112.830 121.215 112.970 ;
        RECT 117.230 112.770 117.550 112.830 ;
        RECT 120.925 112.785 121.215 112.830 ;
        RECT 122.305 112.785 122.595 113.015 ;
        RECT 101.605 112.490 103.200 112.630 ;
        RECT 119.070 112.630 119.390 112.690 ;
        RECT 122.380 112.630 122.520 112.785 ;
        RECT 119.070 112.490 122.520 112.630 ;
        RECT 101.605 112.445 101.895 112.490 ;
        RECT 119.070 112.430 119.390 112.490 ;
        RECT 20.285 112.290 20.575 112.335 ;
        RECT 23.865 112.290 24.155 112.335 ;
        RECT 25.700 112.290 25.990 112.335 ;
        RECT 20.285 112.150 25.990 112.290 ;
        RECT 20.285 112.105 20.575 112.150 ;
        RECT 23.865 112.105 24.155 112.150 ;
        RECT 25.700 112.105 25.990 112.150 ;
        RECT 26.150 112.090 26.470 112.350 ;
        RECT 34.905 112.290 35.195 112.335 ;
        RECT 35.810 112.290 36.130 112.350 ;
        RECT 34.905 112.150 36.130 112.290 ;
        RECT 34.905 112.105 35.195 112.150 ;
        RECT 35.810 112.090 36.130 112.150 ;
        RECT 78.130 112.290 78.450 112.350 ;
        RECT 81.350 112.290 81.670 112.350 ;
        RECT 78.130 112.150 81.670 112.290 ;
        RECT 78.130 112.090 78.450 112.150 ;
        RECT 81.350 112.090 81.670 112.150 ;
        RECT 119.530 112.090 119.850 112.350 ;
        RECT 121.830 112.090 122.150 112.350 ;
        RECT 123.225 112.105 123.515 112.335 ;
        RECT 14.190 111.950 14.510 112.010 ;
        RECT 16.045 111.950 16.335 111.995 ;
        RECT 14.190 111.810 16.335 111.950 ;
        RECT 14.190 111.750 14.510 111.810 ;
        RECT 16.045 111.765 16.335 111.810 ;
        RECT 20.285 111.610 20.575 111.655 ;
        RECT 23.405 111.610 23.695 111.655 ;
        RECT 25.295 111.610 25.585 111.655 ;
        RECT 20.285 111.470 25.585 111.610 ;
        RECT 26.240 111.610 26.380 112.090 ;
        RECT 50.530 111.950 50.850 112.010 ;
        RECT 43.260 111.810 50.850 111.950 ;
        RECT 36.730 111.610 37.050 111.670 ;
        RECT 40.425 111.610 40.715 111.655 ;
        RECT 43.260 111.610 43.400 111.810 ;
        RECT 50.530 111.750 50.850 111.810 ;
        RECT 80.905 111.950 81.195 111.995 ;
        RECT 81.810 111.950 82.130 112.010 ;
        RECT 80.905 111.810 82.130 111.950 ;
        RECT 80.905 111.765 81.195 111.810 ;
        RECT 81.810 111.750 82.130 111.810 ;
        RECT 104.350 111.950 104.670 112.010 ;
        RECT 104.350 111.810 119.760 111.950 ;
        RECT 104.350 111.750 104.670 111.810 ;
        RECT 26.240 111.470 43.400 111.610 ;
        RECT 119.620 111.610 119.760 111.810 ;
        RECT 119.990 111.750 120.310 112.010 ;
        RECT 123.300 111.950 123.440 112.105 ;
        RECT 120.540 111.810 123.440 111.950 ;
        RECT 120.540 111.610 120.680 111.810 ;
        RECT 119.620 111.470 120.680 111.610 ;
        RECT 20.285 111.425 20.575 111.470 ;
        RECT 23.405 111.425 23.695 111.470 ;
        RECT 25.295 111.425 25.585 111.470 ;
        RECT 36.730 111.410 37.050 111.470 ;
        RECT 40.425 111.425 40.715 111.470 ;
        RECT 24.880 111.270 25.170 111.315 ;
        RECT 27.530 111.270 27.850 111.330 ;
        RECT 24.880 111.130 27.850 111.270 ;
        RECT 24.880 111.085 25.170 111.130 ;
        RECT 27.530 111.070 27.850 111.130 ;
        RECT 14.580 110.450 127.740 110.930 ;
        RECT 21.090 110.050 21.410 110.310 ;
        RECT 27.530 110.050 27.850 110.310 ;
        RECT 73.990 110.250 74.310 110.310 ;
        RECT 78.145 110.250 78.435 110.295 ;
        RECT 73.990 110.110 78.435 110.250 ;
        RECT 73.990 110.050 74.310 110.110 ;
        RECT 78.145 110.065 78.435 110.110 ;
        RECT 107.125 109.910 107.415 109.955 ;
        RECT 110.790 109.910 111.110 109.970 ;
        RECT 107.125 109.770 111.110 109.910 ;
        RECT 107.125 109.725 107.415 109.770 ;
        RECT 110.790 109.710 111.110 109.770 ;
        RECT 111.710 109.710 112.030 109.970 ;
        RECT 116.735 109.910 117.025 109.955 ;
        RECT 118.625 109.910 118.915 109.955 ;
        RECT 121.745 109.910 122.035 109.955 ;
        RECT 116.735 109.770 122.035 109.910 ;
        RECT 116.735 109.725 117.025 109.770 ;
        RECT 118.625 109.725 118.915 109.770 ;
        RECT 121.745 109.725 122.035 109.770 ;
        RECT 31.210 109.570 31.530 109.630 ;
        RECT 81.350 109.570 81.670 109.630 ;
        RECT 111.800 109.570 111.940 109.710 ;
        RECT 115.865 109.570 116.155 109.615 ;
        RECT 31.210 109.430 33.280 109.570 ;
        RECT 31.210 109.370 31.530 109.430 ;
        RECT 21.565 109.230 21.855 109.275 ;
        RECT 23.865 109.230 24.155 109.275 ;
        RECT 21.565 109.090 24.155 109.230 ;
        RECT 21.565 109.045 21.855 109.090 ;
        RECT 23.865 109.045 24.155 109.090 ;
        RECT 28.465 109.230 28.755 109.275 ;
        RECT 29.370 109.230 29.690 109.290 ;
        RECT 33.140 109.275 33.280 109.430 ;
        RECT 59.820 109.430 79.740 109.570 ;
        RECT 59.820 109.290 59.960 109.430 ;
        RECT 28.465 109.090 29.690 109.230 ;
        RECT 28.465 109.045 28.755 109.090 ;
        RECT 23.940 108.890 24.080 109.045 ;
        RECT 29.370 109.030 29.690 109.090 ;
        RECT 31.685 109.045 31.975 109.275 ;
        RECT 33.065 109.045 33.355 109.275 ;
        RECT 34.430 109.230 34.750 109.290 ;
        RECT 35.365 109.230 35.655 109.275 ;
        RECT 34.430 109.090 35.655 109.230 ;
        RECT 27.530 108.890 27.850 108.950 ;
        RECT 31.760 108.890 31.900 109.045 ;
        RECT 34.430 109.030 34.750 109.090 ;
        RECT 35.365 109.045 35.655 109.090 ;
        RECT 51.005 109.230 51.295 109.275 ;
        RECT 51.910 109.230 52.230 109.290 ;
        RECT 51.005 109.090 52.230 109.230 ;
        RECT 51.005 109.045 51.295 109.090 ;
        RECT 51.910 109.030 52.230 109.090 ;
        RECT 56.970 109.030 57.290 109.290 ;
        RECT 59.730 109.030 60.050 109.290 ;
        RECT 60.190 109.230 60.510 109.290 ;
        RECT 61.125 109.230 61.415 109.275 ;
        RECT 64.805 109.230 65.095 109.275 ;
        RECT 60.190 109.090 65.095 109.230 ;
        RECT 60.190 109.030 60.510 109.090 ;
        RECT 61.125 109.045 61.415 109.090 ;
        RECT 64.805 109.045 65.095 109.090 ;
        RECT 68.485 109.230 68.775 109.275 ;
        RECT 68.930 109.230 69.250 109.290 ;
        RECT 68.485 109.090 69.250 109.230 ;
        RECT 68.485 109.045 68.775 109.090 ;
        RECT 68.930 109.030 69.250 109.090 ;
        RECT 77.225 109.230 77.515 109.275 ;
        RECT 78.130 109.230 78.450 109.290 ;
        RECT 77.225 109.090 78.450 109.230 ;
        RECT 77.225 109.045 77.515 109.090 ;
        RECT 78.130 109.030 78.450 109.090 ;
        RECT 78.605 109.230 78.895 109.275 ;
        RECT 79.050 109.230 79.370 109.290 ;
        RECT 78.605 109.090 79.370 109.230 ;
        RECT 79.600 109.230 79.740 109.430 ;
        RECT 81.350 109.430 87.560 109.570 ;
        RECT 111.800 109.430 116.155 109.570 ;
        RECT 81.350 109.370 81.670 109.430 ;
        RECT 87.420 109.275 87.560 109.430 ;
        RECT 115.865 109.385 116.155 109.430 ;
        RECT 117.245 109.570 117.535 109.615 ;
        RECT 119.070 109.570 119.390 109.630 ;
        RECT 117.245 109.430 119.390 109.570 ;
        RECT 117.245 109.385 117.535 109.430 ;
        RECT 119.070 109.370 119.390 109.430 ;
        RECT 79.985 109.230 80.275 109.275 ;
        RECT 79.600 109.090 80.275 109.230 ;
        RECT 78.605 109.045 78.895 109.090 ;
        RECT 79.050 109.030 79.370 109.090 ;
        RECT 79.985 109.045 80.275 109.090 ;
        RECT 82.745 109.045 83.035 109.275 ;
        RECT 87.345 109.230 87.635 109.275 ;
        RECT 92.405 109.230 92.695 109.275 ;
        RECT 87.345 109.090 92.695 109.230 ;
        RECT 87.345 109.045 87.635 109.090 ;
        RECT 92.405 109.045 92.695 109.090 ;
        RECT 93.785 109.230 94.075 109.275 ;
        RECT 94.690 109.230 95.010 109.290 ;
        RECT 93.785 109.090 95.010 109.230 ;
        RECT 93.785 109.045 94.075 109.090 ;
        RECT 40.870 108.890 41.190 108.950 ;
        RECT 23.940 108.750 41.190 108.890 ;
        RECT 27.530 108.690 27.850 108.750 ;
        RECT 40.870 108.690 41.190 108.750 ;
        RECT 75.830 108.890 76.150 108.950 ;
        RECT 82.820 108.890 82.960 109.045 ;
        RECT 75.830 108.750 82.960 108.890 ;
        RECT 92.480 108.890 92.620 109.045 ;
        RECT 94.690 109.030 95.010 109.090 ;
        RECT 99.750 109.230 100.070 109.290 ;
        RECT 101.145 109.230 101.435 109.275 ;
        RECT 99.750 109.090 101.435 109.230 ;
        RECT 99.750 109.030 100.070 109.090 ;
        RECT 101.145 109.045 101.435 109.090 ;
        RECT 103.430 109.230 103.750 109.290 ;
        RECT 106.205 109.230 106.495 109.275 ;
        RECT 103.430 109.090 106.495 109.230 ;
        RECT 103.430 109.030 103.750 109.090 ;
        RECT 106.205 109.045 106.495 109.090 ;
        RECT 109.885 109.045 110.175 109.275 ;
        RECT 102.510 108.890 102.830 108.950 ;
        RECT 109.960 108.890 110.100 109.045 ;
        RECT 110.330 109.030 110.650 109.290 ;
        RECT 111.250 109.230 111.570 109.290 ;
        RECT 111.725 109.230 112.015 109.275 ;
        RECT 111.250 109.090 112.015 109.230 ;
        RECT 111.250 109.030 111.570 109.090 ;
        RECT 111.725 109.045 112.015 109.090 ;
        RECT 114.485 109.045 114.775 109.275 ;
        RECT 116.330 109.230 116.620 109.275 ;
        RECT 118.165 109.230 118.455 109.275 ;
        RECT 121.745 109.230 122.035 109.275 ;
        RECT 116.330 109.090 122.035 109.230 ;
        RECT 116.330 109.045 116.620 109.090 ;
        RECT 118.165 109.045 118.455 109.090 ;
        RECT 121.745 109.045 122.035 109.090 ;
        RECT 114.560 108.890 114.700 109.045 ;
        RECT 119.990 108.935 120.310 108.950 ;
        RECT 119.525 108.890 120.310 108.935 ;
        RECT 122.825 108.935 123.115 109.250 ;
        RECT 122.825 108.890 123.415 108.935 ;
        RECT 92.480 108.750 119.300 108.890 ;
        RECT 75.830 108.690 76.150 108.750 ;
        RECT 102.510 108.690 102.830 108.750 ;
        RECT 119.160 108.610 119.300 108.750 ;
        RECT 119.525 108.750 123.415 108.890 ;
        RECT 119.525 108.705 120.310 108.750 ;
        RECT 123.125 108.705 123.415 108.750 ;
        RECT 125.985 108.890 126.275 108.935 ;
        RECT 127.810 108.890 128.130 108.950 ;
        RECT 125.985 108.750 128.130 108.890 ;
        RECT 125.985 108.705 126.275 108.750 ;
        RECT 119.990 108.690 120.310 108.705 ;
        RECT 127.810 108.690 128.130 108.750 ;
        RECT 23.390 108.350 23.710 108.610 ;
        RECT 31.225 108.550 31.515 108.595 ;
        RECT 31.670 108.550 31.990 108.610 ;
        RECT 31.225 108.410 31.990 108.550 ;
        RECT 31.225 108.365 31.515 108.410 ;
        RECT 31.670 108.350 31.990 108.410 ;
        RECT 32.130 108.350 32.450 108.610 ;
        RECT 33.970 108.550 34.290 108.610 ;
        RECT 34.445 108.550 34.735 108.595 ;
        RECT 33.970 108.410 34.735 108.550 ;
        RECT 33.970 108.350 34.290 108.410 ;
        RECT 34.445 108.365 34.735 108.410 ;
        RECT 51.925 108.550 52.215 108.595 ;
        RECT 55.590 108.550 55.910 108.610 ;
        RECT 51.925 108.410 55.910 108.550 ;
        RECT 51.925 108.365 52.215 108.410 ;
        RECT 55.590 108.350 55.910 108.410 ;
        RECT 57.890 108.350 58.210 108.610 ;
        RECT 65.250 108.350 65.570 108.610 ;
        RECT 69.405 108.550 69.695 108.595 ;
        RECT 72.150 108.550 72.470 108.610 ;
        RECT 69.405 108.410 72.470 108.550 ;
        RECT 69.405 108.365 69.695 108.410 ;
        RECT 72.150 108.350 72.470 108.410 ;
        RECT 76.765 108.550 77.055 108.595 ;
        RECT 79.510 108.550 79.830 108.610 ;
        RECT 76.765 108.410 79.830 108.550 ;
        RECT 76.765 108.365 77.055 108.410 ;
        RECT 79.510 108.350 79.830 108.410 ;
        RECT 83.650 108.350 83.970 108.610 ;
        RECT 87.790 108.350 88.110 108.610 ;
        RECT 92.850 108.350 93.170 108.610 ;
        RECT 94.705 108.550 94.995 108.595 ;
        RECT 97.910 108.550 98.230 108.610 ;
        RECT 94.705 108.410 98.230 108.550 ;
        RECT 94.705 108.365 94.995 108.410 ;
        RECT 97.910 108.350 98.230 108.410 ;
        RECT 99.750 108.550 100.070 108.610 ;
        RECT 100.225 108.550 100.515 108.595 ;
        RECT 99.750 108.410 100.515 108.550 ;
        RECT 99.750 108.350 100.070 108.410 ;
        RECT 100.225 108.365 100.515 108.410 ;
        RECT 109.410 108.350 109.730 108.610 ;
        RECT 111.250 108.350 111.570 108.610 ;
        RECT 112.645 108.550 112.935 108.595 ;
        RECT 114.010 108.550 114.330 108.610 ;
        RECT 112.645 108.410 114.330 108.550 ;
        RECT 112.645 108.365 112.935 108.410 ;
        RECT 114.010 108.350 114.330 108.410 ;
        RECT 114.945 108.550 115.235 108.595 ;
        RECT 116.310 108.550 116.630 108.610 ;
        RECT 114.945 108.410 116.630 108.550 ;
        RECT 114.945 108.365 115.235 108.410 ;
        RECT 116.310 108.350 116.630 108.410 ;
        RECT 119.070 108.350 119.390 108.610 ;
        RECT 14.580 107.730 127.740 108.210 ;
        RECT 32.130 107.530 32.450 107.590 ;
        RECT 24.860 107.390 32.450 107.530 ;
        RECT 18.905 107.190 19.195 107.235 ;
        RECT 22.145 107.190 22.795 107.235 ;
        RECT 23.390 107.190 23.710 107.250 ;
        RECT 24.860 107.235 25.000 107.390 ;
        RECT 32.130 107.330 32.450 107.390 ;
        RECT 37.665 107.345 37.955 107.575 ;
        RECT 93.770 107.530 94.090 107.590 ;
        RECT 108.950 107.530 109.270 107.590 ;
        RECT 89.260 107.390 94.090 107.530 ;
        RECT 18.905 107.050 23.710 107.190 ;
        RECT 18.905 107.005 19.495 107.050 ;
        RECT 22.145 107.005 22.795 107.050 ;
        RECT 19.205 106.690 19.495 107.005 ;
        RECT 23.390 106.990 23.710 107.050 ;
        RECT 24.785 107.005 25.075 107.235 ;
        RECT 29.485 107.190 29.775 107.235 ;
        RECT 31.670 107.190 31.990 107.250 ;
        RECT 32.725 107.190 33.375 107.235 ;
        RECT 29.485 107.050 33.375 107.190 ;
        RECT 29.485 107.005 30.075 107.050 ;
        RECT 20.285 106.850 20.575 106.895 ;
        RECT 23.865 106.850 24.155 106.895 ;
        RECT 25.700 106.850 25.990 106.895 ;
        RECT 20.285 106.710 25.990 106.850 ;
        RECT 20.285 106.665 20.575 106.710 ;
        RECT 23.865 106.665 24.155 106.710 ;
        RECT 25.700 106.665 25.990 106.710 ;
        RECT 26.625 106.850 26.915 106.895 ;
        RECT 26.625 106.710 29.600 106.850 ;
        RECT 26.625 106.665 26.915 106.710 ;
        RECT 16.045 106.510 16.335 106.555 ;
        RECT 18.790 106.510 19.110 106.570 ;
        RECT 16.045 106.370 19.110 106.510 ;
        RECT 16.045 106.325 16.335 106.370 ;
        RECT 18.790 106.310 19.110 106.370 ;
        RECT 26.165 106.510 26.455 106.555 ;
        RECT 28.910 106.510 29.230 106.570 ;
        RECT 26.165 106.370 29.230 106.510 ;
        RECT 29.460 106.510 29.600 106.710 ;
        RECT 29.785 106.690 30.075 107.005 ;
        RECT 31.670 106.990 31.990 107.050 ;
        RECT 32.725 107.005 33.375 107.050 ;
        RECT 35.365 107.190 35.655 107.235 ;
        RECT 37.740 107.190 37.880 107.345 ;
        RECT 35.365 107.050 37.880 107.190 ;
        RECT 40.870 107.190 41.190 107.250 ;
        RECT 49.725 107.190 50.015 107.235 ;
        RECT 52.965 107.190 53.615 107.235 ;
        RECT 40.870 107.050 45.240 107.190 ;
        RECT 35.365 107.005 35.655 107.050 ;
        RECT 40.870 106.990 41.190 107.050 ;
        RECT 30.865 106.850 31.155 106.895 ;
        RECT 34.445 106.850 34.735 106.895 ;
        RECT 36.280 106.850 36.570 106.895 ;
        RECT 30.865 106.710 36.570 106.850 ;
        RECT 30.865 106.665 31.155 106.710 ;
        RECT 34.445 106.665 34.735 106.710 ;
        RECT 36.280 106.665 36.570 106.710 ;
        RECT 36.730 106.650 37.050 106.910 ;
        RECT 38.570 106.650 38.890 106.910 ;
        RECT 40.425 106.850 40.715 106.895 ;
        RECT 40.960 106.850 41.100 106.990 ;
        RECT 40.425 106.710 41.100 106.850 ;
        RECT 41.330 106.850 41.650 106.910 ;
        RECT 45.100 106.895 45.240 107.050 ;
        RECT 49.725 107.050 53.615 107.190 ;
        RECT 49.725 107.005 50.315 107.050 ;
        RECT 52.965 107.005 53.615 107.050 ;
        RECT 50.025 106.910 50.315 107.005 ;
        RECT 55.590 106.990 55.910 107.250 ;
        RECT 65.250 107.190 65.570 107.250 ;
        RECT 66.285 107.190 66.575 107.235 ;
        RECT 69.525 107.190 70.175 107.235 ;
        RECT 65.250 107.050 70.175 107.190 ;
        RECT 65.250 106.990 65.570 107.050 ;
        RECT 66.285 107.005 66.875 107.050 ;
        RECT 69.525 107.005 70.175 107.050 ;
        RECT 43.185 106.850 43.475 106.895 ;
        RECT 41.330 106.710 43.475 106.850 ;
        RECT 40.425 106.665 40.715 106.710 ;
        RECT 41.330 106.650 41.650 106.710 ;
        RECT 43.185 106.665 43.475 106.710 ;
        RECT 45.025 106.665 45.315 106.895 ;
        RECT 45.485 106.850 45.775 106.895 ;
        RECT 45.930 106.850 46.250 106.910 ;
        RECT 45.485 106.710 46.250 106.850 ;
        RECT 45.485 106.665 45.775 106.710 ;
        RECT 30.290 106.510 30.610 106.570 ;
        RECT 29.460 106.370 30.610 106.510 ;
        RECT 26.165 106.325 26.455 106.370 ;
        RECT 28.910 106.310 29.230 106.370 ;
        RECT 30.290 106.310 30.610 106.370 ;
        RECT 35.350 106.510 35.670 106.570 ;
        RECT 35.350 106.370 42.480 106.510 ;
        RECT 35.350 106.310 35.670 106.370 ;
        RECT 42.340 106.215 42.480 106.370 ;
        RECT 20.285 106.170 20.575 106.215 ;
        RECT 23.405 106.170 23.695 106.215 ;
        RECT 25.295 106.170 25.585 106.215 ;
        RECT 20.285 106.030 25.585 106.170 ;
        RECT 20.285 105.985 20.575 106.030 ;
        RECT 23.405 105.985 23.695 106.030 ;
        RECT 25.295 105.985 25.585 106.030 ;
        RECT 30.865 106.170 31.155 106.215 ;
        RECT 33.985 106.170 34.275 106.215 ;
        RECT 35.875 106.170 36.165 106.215 ;
        RECT 30.865 106.030 36.165 106.170 ;
        RECT 30.865 105.985 31.155 106.030 ;
        RECT 33.985 105.985 34.275 106.030 ;
        RECT 35.875 105.985 36.165 106.030 ;
        RECT 42.265 105.985 42.555 106.215 ;
        RECT 45.100 106.170 45.240 106.665 ;
        RECT 45.930 106.650 46.250 106.710 ;
        RECT 50.025 106.690 50.390 106.910 ;
        RECT 50.070 106.650 50.390 106.690 ;
        RECT 51.105 106.850 51.395 106.895 ;
        RECT 54.685 106.850 54.975 106.895 ;
        RECT 56.520 106.850 56.810 106.895 ;
        RECT 51.105 106.710 56.810 106.850 ;
        RECT 51.105 106.665 51.395 106.710 ;
        RECT 54.685 106.665 54.975 106.710 ;
        RECT 56.520 106.665 56.810 106.710 ;
        RECT 58.365 106.850 58.655 106.895 ;
        RECT 60.190 106.850 60.510 106.910 ;
        RECT 58.365 106.710 60.510 106.850 ;
        RECT 58.365 106.665 58.655 106.710 ;
        RECT 46.865 106.510 47.155 106.555 ;
        RECT 49.610 106.510 49.930 106.570 ;
        RECT 52.370 106.510 52.690 106.570 ;
        RECT 46.865 106.370 49.930 106.510 ;
        RECT 46.865 106.325 47.155 106.370 ;
        RECT 49.610 106.310 49.930 106.370 ;
        RECT 50.390 106.370 56.740 106.510 ;
        RECT 50.390 106.170 50.530 106.370 ;
        RECT 52.370 106.310 52.690 106.370 ;
        RECT 45.100 106.030 50.530 106.170 ;
        RECT 51.105 106.170 51.395 106.215 ;
        RECT 54.225 106.170 54.515 106.215 ;
        RECT 56.115 106.170 56.405 106.215 ;
        RECT 51.105 106.030 56.405 106.170 ;
        RECT 56.600 106.170 56.740 106.370 ;
        RECT 56.970 106.310 57.290 106.570 ;
        RECT 58.440 106.170 58.580 106.665 ;
        RECT 60.190 106.650 60.510 106.710 ;
        RECT 60.650 106.850 60.970 106.910 ;
        RECT 61.585 106.850 61.875 106.895 ;
        RECT 60.650 106.710 61.875 106.850 ;
        RECT 60.650 106.650 60.970 106.710 ;
        RECT 61.585 106.665 61.875 106.710 ;
        RECT 66.585 106.690 66.875 107.005 ;
        RECT 72.150 106.990 72.470 107.250 ;
        RECT 79.165 107.190 79.455 107.235 ;
        RECT 81.810 107.190 82.130 107.250 ;
        RECT 82.405 107.190 83.055 107.235 ;
        RECT 79.165 107.050 83.055 107.190 ;
        RECT 79.165 107.005 79.755 107.050 ;
        RECT 67.665 106.850 67.955 106.895 ;
        RECT 71.245 106.850 71.535 106.895 ;
        RECT 73.080 106.850 73.370 106.895 ;
        RECT 67.665 106.710 73.370 106.850 ;
        RECT 67.665 106.665 67.955 106.710 ;
        RECT 71.245 106.665 71.535 106.710 ;
        RECT 73.080 106.665 73.370 106.710 ;
        RECT 74.910 106.650 75.230 106.910 ;
        RECT 79.465 106.690 79.755 107.005 ;
        RECT 81.810 106.990 82.130 107.050 ;
        RECT 82.405 107.005 83.055 107.050 ;
        RECT 83.650 107.190 83.970 107.250 ;
        RECT 89.260 107.235 89.400 107.390 ;
        RECT 93.770 107.330 94.090 107.390 ;
        RECT 103.980 107.390 109.270 107.530 ;
        RECT 85.045 107.190 85.335 107.235 ;
        RECT 83.650 107.050 85.335 107.190 ;
        RECT 83.650 106.990 83.970 107.050 ;
        RECT 85.045 107.005 85.335 107.050 ;
        RECT 89.185 107.005 89.475 107.235 ;
        RECT 92.045 107.190 92.335 107.235 ;
        RECT 92.850 107.190 93.170 107.250 ;
        RECT 95.285 107.190 95.935 107.235 ;
        RECT 92.045 107.050 95.935 107.190 ;
        RECT 92.045 107.005 92.635 107.050 ;
        RECT 80.545 106.850 80.835 106.895 ;
        RECT 84.125 106.850 84.415 106.895 ;
        RECT 85.960 106.850 86.250 106.895 ;
        RECT 80.545 106.710 86.250 106.850 ;
        RECT 80.545 106.665 80.835 106.710 ;
        RECT 84.125 106.665 84.415 106.710 ;
        RECT 85.960 106.665 86.250 106.710 ;
        RECT 86.870 106.850 87.190 106.910 ;
        RECT 87.345 106.850 87.635 106.895 ;
        RECT 86.870 106.710 87.635 106.850 ;
        RECT 86.870 106.650 87.190 106.710 ;
        RECT 87.345 106.665 87.635 106.710 ;
        RECT 92.345 106.690 92.635 107.005 ;
        RECT 92.850 106.990 93.170 107.050 ;
        RECT 95.285 107.005 95.935 107.050 ;
        RECT 97.910 106.990 98.230 107.250 ;
        RECT 103.980 107.235 104.120 107.390 ;
        RECT 108.950 107.330 109.270 107.390 ;
        RECT 103.905 107.005 104.195 107.235 ;
        RECT 106.765 107.190 107.055 107.235 ;
        RECT 109.410 107.190 109.730 107.250 ;
        RECT 110.005 107.190 110.655 107.235 ;
        RECT 106.765 107.050 110.655 107.190 ;
        RECT 106.765 107.005 107.355 107.050 ;
        RECT 93.425 106.850 93.715 106.895 ;
        RECT 97.005 106.850 97.295 106.895 ;
        RECT 98.840 106.850 99.130 106.895 ;
        RECT 93.425 106.710 99.130 106.850 ;
        RECT 93.425 106.665 93.715 106.710 ;
        RECT 97.005 106.665 97.295 106.710 ;
        RECT 98.840 106.665 99.130 106.710 ;
        RECT 100.685 106.850 100.975 106.895 ;
        RECT 102.510 106.850 102.830 106.910 ;
        RECT 100.685 106.710 102.830 106.850 ;
        RECT 100.685 106.665 100.975 106.710 ;
        RECT 102.510 106.650 102.830 106.710 ;
        RECT 107.065 106.690 107.355 107.005 ;
        RECT 109.410 106.990 109.730 107.050 ;
        RECT 110.005 107.005 110.655 107.050 ;
        RECT 111.250 107.190 111.570 107.250 ;
        RECT 112.645 107.190 112.935 107.235 ;
        RECT 111.250 107.050 112.935 107.190 ;
        RECT 111.250 106.990 111.570 107.050 ;
        RECT 112.645 107.005 112.935 107.050 ;
        RECT 117.230 106.990 117.550 107.250 ;
        RECT 119.990 107.235 120.310 107.250 ;
        RECT 119.525 107.190 120.310 107.235 ;
        RECT 123.125 107.190 123.415 107.235 ;
        RECT 119.525 107.050 123.415 107.190 ;
        RECT 119.525 107.005 120.310 107.050 ;
        RECT 119.990 106.990 120.310 107.005 ;
        RECT 122.825 107.005 123.415 107.050 ;
        RECT 108.145 106.850 108.435 106.895 ;
        RECT 111.725 106.850 112.015 106.895 ;
        RECT 113.560 106.850 113.850 106.895 ;
        RECT 108.145 106.710 113.850 106.850 ;
        RECT 108.145 106.665 108.435 106.710 ;
        RECT 111.725 106.665 112.015 106.710 ;
        RECT 113.560 106.665 113.850 106.710 ;
        RECT 116.330 106.850 116.620 106.895 ;
        RECT 118.165 106.850 118.455 106.895 ;
        RECT 121.745 106.850 122.035 106.895 ;
        RECT 116.330 106.710 122.035 106.850 ;
        RECT 116.330 106.665 116.620 106.710 ;
        RECT 118.165 106.665 118.455 106.710 ;
        RECT 121.745 106.665 122.035 106.710 ;
        RECT 122.825 106.690 123.115 107.005 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 63.425 106.510 63.715 106.555 ;
        RECT 68.470 106.510 68.790 106.570 ;
        RECT 63.425 106.370 68.790 106.510 ;
        RECT 63.425 106.325 63.715 106.370 ;
        RECT 68.470 106.310 68.790 106.370 ;
        RECT 73.530 106.310 73.850 106.570 ;
        RECT 76.305 106.510 76.595 106.555 ;
        RECT 79.970 106.510 80.290 106.570 ;
        RECT 76.305 106.370 80.290 106.510 ;
        RECT 76.305 106.325 76.595 106.370 ;
        RECT 79.970 106.310 80.290 106.370 ;
        RECT 86.410 106.510 86.730 106.570 ;
        RECT 99.290 106.510 99.610 106.570 ;
        RECT 112.170 106.510 112.490 106.570 ;
        RECT 114.025 106.510 114.315 106.555 ;
        RECT 115.865 106.510 116.155 106.555 ;
        RECT 86.410 106.370 116.155 106.510 ;
        RECT 86.410 106.310 86.730 106.370 ;
        RECT 99.290 106.310 99.610 106.370 ;
        RECT 112.170 106.310 112.490 106.370 ;
        RECT 114.025 106.325 114.315 106.370 ;
        RECT 115.865 106.325 116.155 106.370 ;
        RECT 120.910 106.510 121.230 106.570 ;
        RECT 125.985 106.510 126.275 106.555 ;
        RECT 120.910 106.370 126.275 106.510 ;
        RECT 120.910 106.310 121.230 106.370 ;
        RECT 125.985 106.325 126.275 106.370 ;
        RECT 56.600 106.030 58.580 106.170 ;
        RECT 60.665 106.170 60.955 106.215 ;
        RECT 64.330 106.170 64.650 106.230 ;
        RECT 60.665 106.030 64.650 106.170 ;
        RECT 51.105 105.985 51.395 106.030 ;
        RECT 54.225 105.985 54.515 106.030 ;
        RECT 56.115 105.985 56.405 106.030 ;
        RECT 60.665 105.985 60.955 106.030 ;
        RECT 64.330 105.970 64.650 106.030 ;
        RECT 67.665 106.170 67.955 106.215 ;
        RECT 70.785 106.170 71.075 106.215 ;
        RECT 72.675 106.170 72.965 106.215 ;
        RECT 67.665 106.030 72.965 106.170 ;
        RECT 67.665 105.985 67.955 106.030 ;
        RECT 70.785 105.985 71.075 106.030 ;
        RECT 72.675 105.985 72.965 106.030 ;
        RECT 80.545 106.170 80.835 106.215 ;
        RECT 83.665 106.170 83.955 106.215 ;
        RECT 85.555 106.170 85.845 106.215 ;
        RECT 80.545 106.030 85.845 106.170 ;
        RECT 80.545 105.985 80.835 106.030 ;
        RECT 83.665 105.985 83.955 106.030 ;
        RECT 85.555 105.985 85.845 106.030 ;
        RECT 93.425 106.170 93.715 106.215 ;
        RECT 96.545 106.170 96.835 106.215 ;
        RECT 98.435 106.170 98.725 106.215 ;
        RECT 93.425 106.030 98.725 106.170 ;
        RECT 93.425 105.985 93.715 106.030 ;
        RECT 96.545 105.985 96.835 106.030 ;
        RECT 98.435 105.985 98.725 106.030 ;
        RECT 108.145 106.170 108.435 106.215 ;
        RECT 111.265 106.170 111.555 106.215 ;
        RECT 113.155 106.170 113.445 106.215 ;
        RECT 108.145 106.030 113.445 106.170 ;
        RECT 108.145 105.985 108.435 106.030 ;
        RECT 111.265 105.985 111.555 106.030 ;
        RECT 113.155 105.985 113.445 106.030 ;
        RECT 116.735 106.170 117.025 106.215 ;
        RECT 118.625 106.170 118.915 106.215 ;
        RECT 121.745 106.170 122.035 106.215 ;
        RECT 116.735 106.030 122.035 106.170 ;
        RECT 116.735 105.985 117.025 106.030 ;
        RECT 118.625 105.985 118.915 106.030 ;
        RECT 121.745 105.985 122.035 106.030 ;
        RECT 36.270 105.830 36.590 105.890 ;
        RECT 39.965 105.830 40.255 105.875 ;
        RECT 36.270 105.690 40.255 105.830 ;
        RECT 36.270 105.630 36.590 105.690 ;
        RECT 39.965 105.645 40.255 105.690 ;
        RECT 43.170 105.830 43.490 105.890 ;
        RECT 44.565 105.830 44.855 105.875 ;
        RECT 43.170 105.690 44.855 105.830 ;
        RECT 43.170 105.630 43.490 105.690 ;
        RECT 44.565 105.645 44.855 105.690 ;
        RECT 46.405 105.830 46.695 105.875 ;
        RECT 48.230 105.830 48.550 105.890 ;
        RECT 46.405 105.690 48.550 105.830 ;
        RECT 46.405 105.645 46.695 105.690 ;
        RECT 48.230 105.630 48.550 105.690 ;
        RECT 56.970 105.830 57.290 105.890 ;
        RECT 57.905 105.830 58.195 105.875 ;
        RECT 56.970 105.690 58.195 105.830 ;
        RECT 56.970 105.630 57.290 105.690 ;
        RECT 57.905 105.645 58.195 105.690 ;
        RECT 62.505 105.830 62.795 105.875 ;
        RECT 63.870 105.830 64.190 105.890 ;
        RECT 62.505 105.690 64.190 105.830 ;
        RECT 62.505 105.645 62.795 105.690 ;
        RECT 63.870 105.630 64.190 105.690 ;
        RECT 75.830 105.630 76.150 105.890 ;
        RECT 88.250 105.630 88.570 105.890 ;
        RECT 97.450 105.830 97.770 105.890 ;
        RECT 100.225 105.830 100.515 105.875 ;
        RECT 97.450 105.690 100.515 105.830 ;
        RECT 97.450 105.630 97.770 105.690 ;
        RECT 100.225 105.645 100.515 105.690 ;
        RECT 102.985 105.830 103.275 105.875 ;
        RECT 104.350 105.830 104.670 105.890 ;
        RECT 102.985 105.690 104.670 105.830 ;
        RECT 102.985 105.645 103.275 105.690 ;
        RECT 104.350 105.630 104.670 105.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 14.580 105.010 127.740 105.490 ;
        RECT 28.910 104.810 29.230 104.870 ;
        RECT 36.730 104.810 37.050 104.870 ;
        RECT 28.910 104.670 37.050 104.810 ;
        RECT 28.910 104.610 29.230 104.670 ;
        RECT 36.730 104.610 37.050 104.670 ;
        RECT 50.070 104.810 50.390 104.870 ;
        RECT 51.925 104.810 52.215 104.855 ;
        RECT 50.070 104.670 52.215 104.810 ;
        RECT 50.070 104.610 50.390 104.670 ;
        RECT 51.925 104.625 52.215 104.670 ;
        RECT 56.510 104.810 56.830 104.870 ;
        RECT 73.530 104.810 73.850 104.870 ;
        RECT 56.510 104.670 73.850 104.810 ;
        RECT 56.510 104.610 56.830 104.670 ;
        RECT 29.000 104.175 29.140 104.610 ;
        RECT 29.795 104.470 30.085 104.515 ;
        RECT 31.685 104.470 31.975 104.515 ;
        RECT 34.805 104.470 35.095 104.515 ;
        RECT 29.795 104.330 35.095 104.470 ;
        RECT 29.795 104.285 30.085 104.330 ;
        RECT 31.685 104.285 31.975 104.330 ;
        RECT 34.805 104.285 35.095 104.330 ;
        RECT 43.745 104.470 44.035 104.515 ;
        RECT 46.865 104.470 47.155 104.515 ;
        RECT 48.755 104.470 49.045 104.515 ;
        RECT 50.530 104.470 50.850 104.530 ;
        RECT 56.600 104.470 56.740 104.610 ;
        RECT 43.745 104.330 49.045 104.470 ;
        RECT 43.745 104.285 44.035 104.330 ;
        RECT 46.865 104.285 47.155 104.330 ;
        RECT 48.755 104.285 49.045 104.330 ;
        RECT 50.390 104.330 56.740 104.470 ;
        RECT 57.085 104.470 57.375 104.515 ;
        RECT 60.205 104.470 60.495 104.515 ;
        RECT 62.095 104.470 62.385 104.515 ;
        RECT 57.085 104.330 62.385 104.470 ;
        RECT 50.390 104.270 50.850 104.330 ;
        RECT 57.085 104.285 57.375 104.330 ;
        RECT 60.205 104.285 60.495 104.330 ;
        RECT 62.095 104.285 62.385 104.330 ;
        RECT 28.925 103.945 29.215 104.175 ;
        RECT 30.305 104.130 30.595 104.175 ;
        RECT 35.350 104.130 35.670 104.190 ;
        RECT 36.270 104.130 36.590 104.190 ;
        RECT 30.305 103.990 35.670 104.130 ;
        RECT 30.305 103.945 30.595 103.990 ;
        RECT 35.350 103.930 35.670 103.990 ;
        RECT 35.900 103.990 36.590 104.130 ;
        RECT 27.530 103.590 27.850 103.850 ;
        RECT 29.390 103.790 29.680 103.835 ;
        RECT 31.225 103.790 31.515 103.835 ;
        RECT 34.805 103.790 35.095 103.835 ;
        RECT 35.900 103.810 36.040 103.990 ;
        RECT 36.270 103.930 36.590 103.990 ;
        RECT 48.230 103.930 48.550 104.190 ;
        RECT 49.625 104.130 49.915 104.175 ;
        RECT 50.390 104.130 50.530 104.270 ;
        RECT 49.625 103.990 50.530 104.130 ;
        RECT 57.890 104.130 58.210 104.190 ;
        RECT 63.040 104.175 63.180 104.670 ;
        RECT 73.530 104.610 73.850 104.670 ;
        RECT 79.050 104.810 79.370 104.870 ;
        RECT 125.065 104.810 125.355 104.855 ;
        RECT 79.050 104.670 125.355 104.810 ;
        RECT 79.050 104.610 79.370 104.670 ;
        RECT 125.065 104.625 125.355 104.670 ;
        RECT 67.665 104.470 67.955 104.515 ;
        RECT 70.785 104.470 71.075 104.515 ;
        RECT 72.675 104.470 72.965 104.515 ;
        RECT 67.665 104.330 72.965 104.470 ;
        RECT 67.665 104.285 67.955 104.330 ;
        RECT 70.785 104.285 71.075 104.330 ;
        RECT 72.675 104.285 72.965 104.330 ;
        RECT 80.545 104.470 80.835 104.515 ;
        RECT 83.665 104.470 83.955 104.515 ;
        RECT 85.555 104.470 85.845 104.515 ;
        RECT 80.545 104.330 85.845 104.470 ;
        RECT 80.545 104.285 80.835 104.330 ;
        RECT 83.665 104.285 83.955 104.330 ;
        RECT 85.555 104.285 85.845 104.330 ;
        RECT 91.125 104.470 91.415 104.515 ;
        RECT 94.245 104.470 94.535 104.515 ;
        RECT 96.135 104.470 96.425 104.515 ;
        RECT 91.125 104.330 96.425 104.470 ;
        RECT 91.125 104.285 91.415 104.330 ;
        RECT 94.245 104.285 94.535 104.330 ;
        RECT 96.135 104.285 96.425 104.330 ;
        RECT 106.305 104.470 106.595 104.515 ;
        RECT 109.425 104.470 109.715 104.515 ;
        RECT 111.315 104.470 111.605 104.515 ;
        RECT 106.305 104.330 111.605 104.470 ;
        RECT 106.305 104.285 106.595 104.330 ;
        RECT 109.425 104.285 109.715 104.330 ;
        RECT 111.315 104.285 111.605 104.330 ;
        RECT 113.515 104.470 113.805 104.515 ;
        RECT 115.405 104.470 115.695 104.515 ;
        RECT 118.525 104.470 118.815 104.515 ;
        RECT 113.515 104.330 118.815 104.470 ;
        RECT 113.515 104.285 113.805 104.330 ;
        RECT 115.405 104.285 115.695 104.330 ;
        RECT 118.525 104.285 118.815 104.330 ;
        RECT 61.585 104.130 61.875 104.175 ;
        RECT 57.890 103.990 61.875 104.130 ;
        RECT 49.625 103.945 49.915 103.990 ;
        RECT 57.890 103.930 58.210 103.990 ;
        RECT 61.585 103.945 61.875 103.990 ;
        RECT 62.965 103.945 63.255 104.175 ;
        RECT 63.870 104.130 64.190 104.190 ;
        RECT 72.165 104.130 72.455 104.175 ;
        RECT 63.870 103.990 72.455 104.130 ;
        RECT 63.870 103.930 64.190 103.990 ;
        RECT 72.165 103.945 72.455 103.990 ;
        RECT 73.530 103.930 73.850 104.190 ;
        RECT 75.830 104.130 76.150 104.190 ;
        RECT 85.045 104.130 85.335 104.175 ;
        RECT 75.830 103.990 85.335 104.130 ;
        RECT 75.830 103.930 76.150 103.990 ;
        RECT 85.045 103.945 85.335 103.990 ;
        RECT 86.410 103.930 86.730 104.190 ;
        RECT 88.250 104.130 88.570 104.190 ;
        RECT 95.625 104.130 95.915 104.175 ;
        RECT 88.250 103.990 95.915 104.130 ;
        RECT 88.250 103.930 88.570 103.990 ;
        RECT 95.625 103.945 95.915 103.990 ;
        RECT 97.005 104.130 97.295 104.175 ;
        RECT 99.290 104.130 99.610 104.190 ;
        RECT 97.005 103.990 99.610 104.130 ;
        RECT 97.005 103.945 97.295 103.990 ;
        RECT 99.290 103.930 99.610 103.990 ;
        RECT 110.790 103.930 111.110 104.190 ;
        RECT 112.170 104.130 112.490 104.190 ;
        RECT 112.645 104.130 112.935 104.175 ;
        RECT 112.170 103.990 112.935 104.130 ;
        RECT 112.170 103.930 112.490 103.990 ;
        RECT 112.645 103.945 112.935 103.990 ;
        RECT 114.010 103.930 114.330 104.190 ;
        RECT 115.850 104.130 116.170 104.190 ;
        RECT 122.765 104.130 123.055 104.175 ;
        RECT 115.850 103.990 123.055 104.130 ;
        RECT 115.850 103.930 116.170 103.990 ;
        RECT 122.765 103.945 123.055 103.990 ;
        RECT 29.390 103.650 35.095 103.790 ;
        RECT 29.390 103.605 29.680 103.650 ;
        RECT 31.225 103.605 31.515 103.650 ;
        RECT 34.805 103.605 35.095 103.650 ;
        RECT 35.885 103.495 36.175 103.810 ;
        RECT 32.585 103.450 33.235 103.495 ;
        RECT 35.885 103.450 36.475 103.495 ;
        RECT 32.585 103.310 36.475 103.450 ;
        RECT 32.585 103.265 33.235 103.310 ;
        RECT 36.185 103.265 36.475 103.310 ;
        RECT 39.030 103.250 39.350 103.510 ;
        RECT 42.665 103.495 42.955 103.810 ;
        RECT 43.745 103.790 44.035 103.835 ;
        RECT 47.325 103.790 47.615 103.835 ;
        RECT 49.160 103.790 49.450 103.835 ;
        RECT 43.745 103.650 49.450 103.790 ;
        RECT 43.745 103.605 44.035 103.650 ;
        RECT 47.325 103.605 47.615 103.650 ;
        RECT 49.160 103.605 49.450 103.650 ;
        RECT 52.370 103.590 52.690 103.850 ;
        RECT 39.505 103.265 39.795 103.495 ;
        RECT 42.365 103.450 42.955 103.495 ;
        RECT 43.170 103.450 43.490 103.510 ;
        RECT 45.605 103.450 46.255 103.495 ;
        RECT 42.365 103.310 46.255 103.450 ;
        RECT 42.365 103.265 42.655 103.310 ;
        RECT 27.990 102.910 28.310 103.170 ;
        RECT 39.580 103.110 39.720 103.265 ;
        RECT 43.170 103.250 43.490 103.310 ;
        RECT 45.605 103.265 46.255 103.310 ;
        RECT 52.845 103.450 53.135 103.495 ;
        RECT 54.670 103.450 54.990 103.510 ;
        RECT 56.005 103.495 56.295 103.810 ;
        RECT 57.085 103.790 57.375 103.835 ;
        RECT 60.665 103.790 60.955 103.835 ;
        RECT 62.500 103.790 62.790 103.835 ;
        RECT 57.085 103.650 62.790 103.790 ;
        RECT 57.085 103.605 57.375 103.650 ;
        RECT 60.665 103.605 60.955 103.650 ;
        RECT 62.500 103.605 62.790 103.650 ;
        RECT 52.845 103.310 54.990 103.450 ;
        RECT 52.845 103.265 53.135 103.310 ;
        RECT 54.670 103.250 54.990 103.310 ;
        RECT 55.705 103.450 56.295 103.495 ;
        RECT 56.510 103.450 56.830 103.510 ;
        RECT 58.945 103.450 59.595 103.495 ;
        RECT 55.705 103.310 59.595 103.450 ;
        RECT 55.705 103.265 55.995 103.310 ;
        RECT 56.510 103.250 56.830 103.310 ;
        RECT 58.945 103.265 59.595 103.310 ;
        RECT 61.110 103.450 61.430 103.510 ;
        RECT 63.425 103.450 63.715 103.495 ;
        RECT 61.110 103.310 63.715 103.450 ;
        RECT 61.110 103.250 61.430 103.310 ;
        RECT 63.425 103.265 63.715 103.310 ;
        RECT 64.330 103.450 64.650 103.510 ;
        RECT 66.585 103.495 66.875 103.810 ;
        RECT 67.665 103.790 67.955 103.835 ;
        RECT 71.245 103.790 71.535 103.835 ;
        RECT 73.080 103.790 73.370 103.835 ;
        RECT 79.510 103.810 79.830 103.850 ;
        RECT 67.665 103.650 73.370 103.790 ;
        RECT 67.665 103.605 67.955 103.650 ;
        RECT 71.245 103.605 71.535 103.650 ;
        RECT 73.080 103.605 73.370 103.650 ;
        RECT 79.465 103.590 79.830 103.810 ;
        RECT 80.545 103.790 80.835 103.835 ;
        RECT 84.125 103.790 84.415 103.835 ;
        RECT 85.960 103.790 86.250 103.835 ;
        RECT 80.545 103.650 86.250 103.790 ;
        RECT 80.545 103.605 80.835 103.650 ;
        RECT 84.125 103.605 84.415 103.650 ;
        RECT 85.960 103.605 86.250 103.650 ;
        RECT 66.285 103.450 66.875 103.495 ;
        RECT 69.525 103.450 70.175 103.495 ;
        RECT 64.330 103.310 70.175 103.450 ;
        RECT 64.330 103.250 64.650 103.310 ;
        RECT 66.285 103.265 66.575 103.310 ;
        RECT 69.525 103.265 70.175 103.310 ;
        RECT 73.990 103.450 74.310 103.510 ;
        RECT 79.465 103.495 79.755 103.590 ;
        RECT 76.305 103.450 76.595 103.495 ;
        RECT 73.990 103.310 76.595 103.450 ;
        RECT 73.990 103.250 74.310 103.310 ;
        RECT 76.305 103.265 76.595 103.310 ;
        RECT 79.165 103.450 79.755 103.495 ;
        RECT 82.405 103.450 83.055 103.495 ;
        RECT 79.165 103.310 83.055 103.450 ;
        RECT 79.165 103.265 79.455 103.310 ;
        RECT 82.405 103.265 83.055 103.310 ;
        RECT 86.870 103.250 87.190 103.510 ;
        RECT 87.790 103.450 88.110 103.510 ;
        RECT 90.045 103.495 90.335 103.810 ;
        RECT 91.125 103.790 91.415 103.835 ;
        RECT 94.705 103.790 94.995 103.835 ;
        RECT 96.540 103.790 96.830 103.835 ;
        RECT 91.125 103.650 96.830 103.790 ;
        RECT 91.125 103.605 91.415 103.650 ;
        RECT 94.705 103.605 94.995 103.650 ;
        RECT 96.540 103.605 96.830 103.650 ;
        RECT 89.745 103.450 90.335 103.495 ;
        RECT 92.985 103.450 93.635 103.495 ;
        RECT 87.790 103.310 93.635 103.450 ;
        RECT 87.790 103.250 88.110 103.310 ;
        RECT 89.745 103.265 90.035 103.310 ;
        RECT 92.985 103.265 93.635 103.310 ;
        RECT 102.065 103.450 102.355 103.495 ;
        RECT 103.890 103.450 104.210 103.510 ;
        RECT 102.065 103.310 104.210 103.450 ;
        RECT 102.065 103.265 102.355 103.310 ;
        RECT 103.890 103.250 104.210 103.310 ;
        RECT 104.350 103.450 104.670 103.510 ;
        RECT 105.225 103.495 105.515 103.810 ;
        RECT 106.305 103.790 106.595 103.835 ;
        RECT 109.885 103.790 110.175 103.835 ;
        RECT 111.720 103.790 112.010 103.835 ;
        RECT 106.305 103.650 112.010 103.790 ;
        RECT 106.305 103.605 106.595 103.650 ;
        RECT 109.885 103.605 110.175 103.650 ;
        RECT 111.720 103.605 112.010 103.650 ;
        RECT 113.110 103.790 113.400 103.835 ;
        RECT 114.945 103.790 115.235 103.835 ;
        RECT 118.525 103.790 118.815 103.835 ;
        RECT 113.110 103.650 118.815 103.790 ;
        RECT 113.110 103.605 113.400 103.650 ;
        RECT 114.945 103.605 115.235 103.650 ;
        RECT 118.525 103.605 118.815 103.650 ;
        RECT 116.310 103.495 116.630 103.510 ;
        RECT 119.605 103.495 119.895 103.810 ;
        RECT 125.970 103.590 126.290 103.850 ;
        RECT 104.925 103.450 105.515 103.495 ;
        RECT 108.165 103.450 108.815 103.495 ;
        RECT 104.350 103.310 108.815 103.450 ;
        RECT 104.350 103.250 104.670 103.310 ;
        RECT 104.925 103.265 105.215 103.310 ;
        RECT 108.165 103.265 108.815 103.310 ;
        RECT 116.305 103.450 116.955 103.495 ;
        RECT 119.605 103.450 120.195 103.495 ;
        RECT 116.305 103.310 120.195 103.450 ;
        RECT 116.305 103.265 116.955 103.310 ;
        RECT 119.905 103.265 120.195 103.310 ;
        RECT 116.310 103.250 116.630 103.265 ;
        RECT 44.090 103.110 44.410 103.170 ;
        RECT 39.580 102.970 44.410 103.110 ;
        RECT 44.090 102.910 44.410 102.970 ;
        RECT 14.580 102.290 127.740 102.770 ;
        RECT 119.990 101.890 120.310 102.150 ;
        RECT 27.645 101.750 27.935 101.795 ;
        RECT 30.885 101.750 31.535 101.795 ;
        RECT 27.645 101.610 31.535 101.750 ;
        RECT 27.645 101.565 28.235 101.610 ;
        RECT 30.885 101.565 31.535 101.610 ;
        RECT 33.525 101.750 33.815 101.795 ;
        RECT 33.970 101.750 34.290 101.810 ;
        RECT 97.450 101.795 97.770 101.810 ;
        RECT 33.525 101.610 34.290 101.750 ;
        RECT 33.525 101.565 33.815 101.610 ;
        RECT 27.945 101.470 28.235 101.565 ;
        RECT 33.970 101.550 34.290 101.610 ;
        RECT 93.885 101.750 94.175 101.795 ;
        RECT 97.125 101.750 97.775 101.795 ;
        RECT 93.885 101.610 97.775 101.750 ;
        RECT 93.885 101.565 94.475 101.610 ;
        RECT 97.125 101.565 97.775 101.610 ;
        RECT 27.945 101.250 28.310 101.470 ;
        RECT 27.990 101.210 28.310 101.250 ;
        RECT 29.025 101.410 29.315 101.455 ;
        RECT 32.605 101.410 32.895 101.455 ;
        RECT 34.440 101.410 34.730 101.455 ;
        RECT 29.025 101.270 34.730 101.410 ;
        RECT 29.025 101.225 29.315 101.270 ;
        RECT 32.605 101.225 32.895 101.270 ;
        RECT 34.440 101.225 34.730 101.270 ;
        RECT 34.905 101.410 35.195 101.455 ;
        RECT 36.730 101.410 37.050 101.470 ;
        RECT 34.905 101.270 37.050 101.410 ;
        RECT 34.905 101.225 35.195 101.270 ;
        RECT 36.730 101.210 37.050 101.270 ;
        RECT 94.185 101.250 94.475 101.565 ;
        RECT 97.450 101.550 97.770 101.565 ;
        RECT 99.750 101.550 100.070 101.810 ;
        RECT 95.265 101.410 95.555 101.455 ;
        RECT 98.845 101.410 99.135 101.455 ;
        RECT 100.680 101.410 100.970 101.455 ;
        RECT 95.265 101.270 100.970 101.410 ;
        RECT 95.265 101.225 95.555 101.270 ;
        RECT 98.845 101.225 99.135 101.270 ;
        RECT 100.680 101.225 100.970 101.270 ;
        RECT 119.530 101.210 119.850 101.470 ;
        RECT 24.785 101.070 25.075 101.115 ;
        RECT 26.150 101.070 26.470 101.130 ;
        RECT 24.785 100.930 26.470 101.070 ;
        RECT 24.785 100.885 25.075 100.930 ;
        RECT 26.150 100.870 26.470 100.930 ;
        RECT 91.025 101.070 91.315 101.115 ;
        RECT 97.910 101.070 98.230 101.130 ;
        RECT 91.025 100.930 98.230 101.070 ;
        RECT 91.025 100.885 91.315 100.930 ;
        RECT 97.910 100.870 98.230 100.930 ;
        RECT 99.290 101.070 99.610 101.130 ;
        RECT 101.145 101.070 101.435 101.115 ;
        RECT 99.290 100.930 101.435 101.070 ;
        RECT 99.290 100.870 99.610 100.930 ;
        RECT 101.145 100.885 101.435 100.930 ;
        RECT 29.025 100.730 29.315 100.775 ;
        RECT 32.145 100.730 32.435 100.775 ;
        RECT 34.035 100.730 34.325 100.775 ;
        RECT 29.025 100.590 34.325 100.730 ;
        RECT 29.025 100.545 29.315 100.590 ;
        RECT 32.145 100.545 32.435 100.590 ;
        RECT 34.035 100.545 34.325 100.590 ;
        RECT 95.265 100.730 95.555 100.775 ;
        RECT 98.385 100.730 98.675 100.775 ;
        RECT 100.275 100.730 100.565 100.775 ;
        RECT 95.265 100.590 100.565 100.730 ;
        RECT 95.265 100.545 95.555 100.590 ;
        RECT 98.385 100.545 98.675 100.590 ;
        RECT 100.275 100.545 100.565 100.590 ;
        RECT 14.580 99.570 127.740 100.050 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 16.800 211.145 18.680 211.515 ;
        RECT 46.800 211.145 48.680 211.515 ;
        RECT 76.800 211.145 78.680 211.515 ;
        RECT 106.800 211.145 108.680 211.515 ;
        RECT 31.800 208.425 33.680 208.795 ;
        RECT 61.800 208.425 63.680 208.795 ;
        RECT 91.800 208.425 93.680 208.795 ;
        RECT 121.800 208.425 123.680 208.795 ;
        RECT 73.560 207.600 73.820 207.920 ;
        RECT 66.200 206.920 66.460 207.240 ;
        RECT 73.100 206.920 73.360 207.240 ;
        RECT 16.800 205.705 18.680 206.075 ;
        RECT 46.800 205.705 48.680 206.075 ;
        RECT 66.260 204.860 66.400 206.920 ;
        RECT 66.200 204.540 66.460 204.860 ;
        RECT 63.900 204.200 64.160 204.520 ;
        RECT 31.800 202.985 33.680 203.355 ;
        RECT 61.800 202.985 63.680 203.355 ;
        RECT 63.960 202.820 64.100 204.200 ;
        RECT 64.820 203.520 65.080 203.840 ;
        RECT 63.900 202.500 64.160 202.820 ;
        RECT 61.140 201.820 61.400 202.140 ;
        RECT 16.800 200.265 18.680 200.635 ;
        RECT 46.800 200.265 48.680 200.635 ;
        RECT 61.200 200.100 61.340 201.820 ;
        RECT 61.140 199.780 61.400 200.100 ;
        RECT 31.800 197.545 33.680 197.915 ;
        RECT 61.800 197.545 63.680 197.915 ;
        RECT 50.560 196.380 50.820 196.700 ;
        RECT 49.180 196.040 49.440 196.360 ;
        RECT 16.800 194.825 18.680 195.195 ;
        RECT 46.800 194.825 48.680 195.195 ;
        RECT 49.240 194.320 49.380 196.040 ;
        RECT 50.620 194.660 50.760 196.380 ;
        RECT 53.320 195.360 53.580 195.680 ;
        RECT 57.920 195.360 58.180 195.680 ;
        RECT 50.560 194.570 50.820 194.660 ;
        RECT 49.700 194.430 50.820 194.570 ;
        RECT 49.180 194.000 49.440 194.320 ;
        RECT 45.960 193.660 46.220 193.980 ;
        RECT 31.800 192.105 33.680 192.475 ;
        RECT 41.360 190.940 41.620 191.260 ;
        RECT 39.060 190.260 39.320 190.580 ;
        RECT 16.800 189.385 18.680 189.755 ;
        RECT 28.480 187.880 28.740 188.200 ;
        RECT 36.300 187.880 36.560 188.200 ;
        RECT 22.960 185.500 23.220 185.820 ;
        RECT 16.800 183.945 18.680 184.315 ;
        RECT 23.020 183.780 23.160 185.500 ;
        RECT 28.540 185.140 28.680 187.880 ;
        RECT 31.800 186.665 33.680 187.035 ;
        RECT 36.360 185.480 36.500 187.880 ;
        RECT 37.680 187.200 37.940 187.520 ;
        RECT 36.300 185.160 36.560 185.480 ;
        RECT 28.480 184.820 28.740 185.140 ;
        RECT 29.860 184.480 30.120 184.800 ;
        RECT 30.320 184.480 30.580 184.800 ;
        RECT 22.960 183.460 23.220 183.780 ;
        RECT 29.920 183.100 30.060 184.480 ;
        RECT 30.380 183.780 30.520 184.480 ;
        RECT 30.320 183.460 30.580 183.780 ;
        RECT 34.000 183.120 34.260 183.440 ;
        RECT 29.860 182.780 30.120 183.100 ;
        RECT 31.800 181.225 33.680 181.595 ;
        RECT 34.060 179.700 34.200 183.120 ;
        RECT 35.840 182.780 36.100 183.100 ;
        RECT 26.180 179.380 26.440 179.700 ;
        RECT 27.560 179.380 27.820 179.700 ;
        RECT 34.000 179.380 34.260 179.700 ;
        RECT 34.920 179.380 35.180 179.700 ;
        RECT 16.800 178.505 18.680 178.875 ;
        RECT 26.240 175.620 26.380 179.380 ;
        RECT 27.620 178.340 27.760 179.380 ;
        RECT 27.560 178.020 27.820 178.340 ;
        RECT 30.320 177.000 30.580 177.320 ;
        RECT 28.020 176.320 28.280 176.640 ;
        RECT 26.180 175.300 26.440 175.620 ;
        RECT 28.080 174.260 28.220 176.320 ;
        RECT 28.020 173.940 28.280 174.260 ;
        RECT 16.800 173.065 18.680 173.435 ;
        RECT 30.380 169.160 30.520 177.000 ;
        RECT 31.800 175.785 33.680 176.155 ;
        RECT 34.060 174.260 34.200 179.380 ;
        RECT 34.460 176.320 34.720 176.640 ;
        RECT 34.520 174.600 34.660 176.320 ;
        RECT 34.460 174.280 34.720 174.600 ;
        RECT 34.000 173.940 34.260 174.260 ;
        RECT 31.800 170.345 33.680 170.715 ;
        RECT 30.320 168.840 30.580 169.160 ;
        RECT 29.860 168.160 30.120 168.480 ;
        RECT 34.000 168.160 34.260 168.480 ;
        RECT 16.800 167.625 18.680 167.995 ;
        RECT 29.920 167.120 30.060 168.160 ;
        RECT 24.800 166.800 25.060 167.120 ;
        RECT 29.860 166.800 30.120 167.120 ;
        RECT 24.860 164.740 25.000 166.800 ;
        RECT 27.100 166.120 27.360 166.440 ;
        RECT 24.800 164.420 25.060 164.740 ;
        RECT 27.160 163.720 27.300 166.120 ;
        RECT 29.860 165.780 30.120 166.100 ;
        RECT 28.480 165.440 28.740 165.760 ;
        RECT 28.540 164.060 28.680 165.440 ;
        RECT 28.480 163.740 28.740 164.060 ;
        RECT 28.940 163.740 29.200 164.060 ;
        RECT 26.640 163.400 26.900 163.720 ;
        RECT 27.100 163.400 27.360 163.720 ;
        RECT 16.800 162.185 18.680 162.555 ;
        RECT 26.700 162.020 26.840 163.400 ;
        RECT 29.000 163.380 29.140 163.740 ;
        RECT 28.940 163.060 29.200 163.380 ;
        RECT 26.640 161.700 26.900 162.020 ;
        RECT 18.820 161.360 19.080 161.680 ;
        RECT 18.880 159.300 19.020 161.360 ;
        RECT 29.000 161.340 29.140 163.060 ;
        RECT 29.920 162.020 30.060 165.780 ;
        RECT 31.800 164.905 33.680 165.275 ;
        RECT 34.060 163.720 34.200 168.160 ;
        RECT 34.460 166.460 34.720 166.780 ;
        RECT 34.000 163.400 34.260 163.720 ;
        RECT 34.520 162.020 34.660 166.460 ;
        RECT 29.860 161.700 30.120 162.020 ;
        RECT 34.460 161.700 34.720 162.020 ;
        RECT 31.240 161.360 31.500 161.680 ;
        RECT 34.980 161.420 35.120 179.380 ;
        RECT 35.380 177.000 35.640 177.320 ;
        RECT 35.440 172.900 35.580 177.000 ;
        RECT 35.380 172.580 35.640 172.900 ;
        RECT 35.900 171.880 36.040 182.780 ;
        RECT 35.840 171.560 36.100 171.880 ;
        RECT 35.380 170.880 35.640 171.200 ;
        RECT 36.360 170.940 36.500 185.160 ;
        RECT 37.740 185.140 37.880 187.200 ;
        RECT 39.120 186.500 39.260 190.260 ;
        RECT 39.060 186.180 39.320 186.500 ;
        RECT 41.420 185.820 41.560 190.940 ;
        RECT 45.040 190.600 45.300 190.920 ;
        RECT 44.580 187.880 44.840 188.200 ;
        RECT 44.640 186.160 44.780 187.880 ;
        RECT 44.580 185.840 44.840 186.160 ;
        RECT 38.140 185.500 38.400 185.820 ;
        RECT 41.360 185.500 41.620 185.820 ;
        RECT 37.680 184.820 37.940 185.140 ;
        RECT 37.740 183.100 37.880 184.820 ;
        RECT 37.680 182.780 37.940 183.100 ;
        RECT 37.220 179.720 37.480 180.040 ;
        RECT 36.760 179.040 37.020 179.360 ;
        RECT 36.820 177.320 36.960 179.040 ;
        RECT 36.760 177.000 37.020 177.320 ;
        RECT 27.100 161.020 27.360 161.340 ;
        RECT 28.940 161.020 29.200 161.340 ;
        RECT 25.720 160.680 25.980 161.000 ;
        RECT 21.580 160.000 21.840 160.320 ;
        RECT 18.820 158.980 19.080 159.300 ;
        RECT 21.640 158.620 21.780 160.000 ;
        RECT 25.780 159.300 25.920 160.680 ;
        RECT 25.720 158.980 25.980 159.300 ;
        RECT 21.120 158.300 21.380 158.620 ;
        RECT 21.580 158.300 21.840 158.620 ;
        RECT 19.280 157.280 19.540 157.600 ;
        RECT 16.800 156.745 18.680 157.115 ;
        RECT 19.340 156.240 19.480 157.280 ;
        RECT 19.280 155.920 19.540 156.240 ;
        RECT 21.180 153.180 21.320 158.300 ;
        RECT 22.040 157.280 22.300 157.600 ;
        RECT 22.100 156.580 22.240 157.280 ;
        RECT 22.040 156.260 22.300 156.580 ;
        RECT 22.100 153.180 22.240 156.260 ;
        RECT 27.160 155.900 27.300 161.020 ;
        RECT 30.780 160.680 31.040 161.000 ;
        RECT 30.840 158.960 30.980 160.680 ;
        RECT 31.300 159.300 31.440 161.360 ;
        RECT 34.000 161.020 34.260 161.340 ;
        RECT 34.520 161.280 35.120 161.420 ;
        RECT 34.060 160.320 34.200 161.020 ;
        RECT 34.000 160.000 34.260 160.320 ;
        RECT 31.800 159.465 33.680 159.835 ;
        RECT 31.240 158.980 31.500 159.300 ;
        RECT 30.780 158.640 31.040 158.960 ;
        RECT 29.860 158.300 30.120 158.620 ;
        RECT 27.100 155.580 27.360 155.900 ;
        RECT 27.560 155.580 27.820 155.900 ;
        RECT 27.620 153.860 27.760 155.580 ;
        RECT 27.560 153.540 27.820 153.860 ;
        RECT 21.120 152.860 21.380 153.180 ;
        RECT 22.040 152.860 22.300 153.180 ;
        RECT 16.800 151.305 18.680 151.675 ;
        RECT 20.200 150.480 20.460 150.800 ;
        RECT 16.800 145.865 18.680 146.235 ;
        RECT 20.260 145.700 20.400 150.480 ;
        RECT 21.180 147.740 21.320 152.860 ;
        RECT 22.500 151.840 22.760 152.160 ;
        RECT 22.560 150.120 22.700 151.840 ;
        RECT 29.920 150.460 30.060 158.300 ;
        RECT 30.840 155.560 30.980 158.640 ;
        RECT 32.160 157.960 32.420 158.280 ;
        RECT 31.240 155.580 31.500 155.900 ;
        RECT 30.780 155.240 31.040 155.560 ;
        RECT 31.300 152.160 31.440 155.580 ;
        RECT 32.220 155.220 32.360 157.960 ;
        RECT 33.540 156.260 33.800 156.580 ;
        RECT 33.600 155.900 33.740 156.260 ;
        RECT 33.540 155.580 33.800 155.900 ;
        RECT 34.000 155.240 34.260 155.560 ;
        RECT 32.160 154.900 32.420 155.220 ;
        RECT 31.800 154.025 33.680 154.395 ;
        RECT 33.540 152.180 33.800 152.500 ;
        RECT 31.240 151.840 31.500 152.160 ;
        RECT 31.300 150.800 31.440 151.840 ;
        RECT 33.600 151.140 33.740 152.180 ;
        RECT 33.540 150.820 33.800 151.140 ;
        RECT 31.240 150.480 31.500 150.800 ;
        RECT 29.860 150.140 30.120 150.460 ;
        RECT 22.500 149.800 22.760 150.120 ;
        RECT 24.800 149.800 25.060 150.120 ;
        RECT 21.120 147.420 21.380 147.740 ;
        RECT 22.560 146.720 22.700 149.800 ;
        RECT 24.860 148.420 25.000 149.800 ;
        RECT 24.800 148.100 25.060 148.420 ;
        RECT 28.480 147.760 28.740 148.080 ;
        RECT 22.960 146.740 23.220 147.060 ;
        RECT 22.500 146.400 22.760 146.720 ;
        RECT 23.020 145.700 23.160 146.740 ;
        RECT 28.540 146.720 28.680 147.760 ;
        RECT 28.480 146.400 28.740 146.720 ;
        RECT 28.940 146.400 29.200 146.720 ;
        RECT 20.200 145.380 20.460 145.700 ;
        RECT 22.960 145.380 23.220 145.700 ;
        RECT 29.000 144.680 29.140 146.400 ;
        RECT 29.920 145.100 30.060 150.140 ;
        RECT 31.300 147.400 31.440 150.480 ;
        RECT 31.800 148.585 33.680 148.955 ;
        RECT 34.060 147.740 34.200 155.240 ;
        RECT 34.000 147.420 34.260 147.740 ;
        RECT 31.240 147.080 31.500 147.400 ;
        RECT 29.920 145.020 30.520 145.100 ;
        RECT 29.920 144.960 30.580 145.020 ;
        RECT 28.940 144.360 29.200 144.680 ;
        RECT 29.920 144.000 30.060 144.960 ;
        RECT 30.320 144.700 30.580 144.960 ;
        RECT 29.860 143.680 30.120 144.000 ;
        RECT 31.800 143.145 33.680 143.515 ;
        RECT 34.520 142.300 34.660 161.280 ;
        RECT 34.920 160.000 35.180 160.320 ;
        RECT 34.980 157.600 35.120 160.000 ;
        RECT 34.920 157.280 35.180 157.600 ;
        RECT 34.980 156.580 35.120 157.280 ;
        RECT 34.920 156.260 35.180 156.580 ;
        RECT 34.920 151.840 35.180 152.160 ;
        RECT 34.460 141.980 34.720 142.300 ;
        RECT 34.980 141.960 35.120 151.840 ;
        RECT 34.920 141.640 35.180 141.960 ;
        RECT 29.400 140.960 29.660 141.280 ;
        RECT 16.800 140.425 18.680 140.795 ;
        RECT 19.280 139.600 19.540 139.920 ;
        RECT 18.820 135.520 19.080 135.840 ;
        RECT 16.800 134.985 18.680 135.355 ;
        RECT 18.880 134.140 19.020 135.520 ;
        RECT 19.340 134.820 19.480 139.600 ;
        RECT 23.420 138.920 23.680 139.240 ;
        RECT 22.500 138.240 22.760 138.560 ;
        RECT 21.580 136.540 21.840 136.860 ;
        RECT 19.280 134.500 19.540 134.820 ;
        RECT 21.640 134.220 21.780 136.540 ;
        RECT 22.560 136.520 22.700 138.240 ;
        RECT 22.500 136.200 22.760 136.520 ;
        RECT 22.040 135.520 22.300 135.840 ;
        RECT 22.100 134.820 22.240 135.520 ;
        RECT 22.040 134.500 22.300 134.820 ;
        RECT 18.820 133.820 19.080 134.140 ;
        RECT 21.640 134.080 22.240 134.220 ;
        RECT 22.100 133.800 22.240 134.080 ;
        RECT 19.740 133.480 20.000 133.800 ;
        RECT 22.040 133.480 22.300 133.800 ;
        RECT 16.800 129.545 18.680 129.915 ;
        RECT 19.800 125.980 19.940 133.480 ;
        RECT 22.100 131.420 22.240 133.480 ;
        RECT 22.040 131.100 22.300 131.420 ;
        RECT 21.120 128.720 21.380 129.040 ;
        RECT 19.740 125.660 20.000 125.980 ;
        RECT 16.800 124.105 18.680 124.475 ;
        RECT 16.800 118.665 18.680 119.035 ;
        RECT 19.800 117.900 19.940 125.660 ;
        RECT 21.180 125.640 21.320 128.720 ;
        RECT 21.120 125.320 21.380 125.640 ;
        RECT 22.100 122.920 22.240 131.100 ;
        RECT 22.560 130.400 22.700 136.200 ;
        RECT 23.480 133.460 23.620 138.920 ;
        RECT 28.480 135.520 28.740 135.840 ;
        RECT 23.420 133.140 23.680 133.460 ;
        RECT 28.540 131.080 28.680 135.520 ;
        RECT 28.940 133.480 29.200 133.800 ;
        RECT 29.000 132.100 29.140 133.480 ;
        RECT 28.940 131.780 29.200 132.100 ;
        RECT 28.480 130.760 28.740 131.080 ;
        RECT 23.420 130.420 23.680 130.740 ;
        RECT 22.500 130.080 22.760 130.400 ;
        RECT 22.960 130.080 23.220 130.400 ;
        RECT 22.560 127.680 22.700 130.080 ;
        RECT 22.500 127.360 22.760 127.680 ;
        RECT 23.020 125.640 23.160 130.080 ;
        RECT 23.480 129.380 23.620 130.420 ;
        RECT 23.420 129.060 23.680 129.380 ;
        RECT 22.960 125.320 23.220 125.640 ;
        RECT 23.480 123.940 23.620 129.060 ;
        RECT 23.880 128.040 24.140 128.360 ;
        RECT 23.940 126.660 24.080 128.040 ;
        RECT 23.880 126.340 24.140 126.660 ;
        RECT 22.500 123.620 22.760 123.940 ;
        RECT 23.420 123.620 23.680 123.940 ;
        RECT 22.040 122.600 22.300 122.920 ;
        RECT 22.100 120.880 22.240 122.600 ;
        RECT 22.040 120.560 22.300 120.880 ;
        RECT 22.560 120.540 22.700 123.620 ;
        RECT 26.640 121.920 26.900 122.240 ;
        RECT 22.500 120.220 22.760 120.540 ;
        RECT 21.120 119.200 21.380 119.520 ;
        RECT 19.340 117.820 19.940 117.900 ;
        RECT 19.280 117.760 19.940 117.820 ;
        RECT 19.280 117.500 19.540 117.760 ;
        RECT 19.800 115.100 19.940 117.760 ;
        RECT 19.740 114.780 20.000 115.100 ;
        RECT 21.180 114.760 21.320 119.200 ;
        RECT 22.560 118.500 22.700 120.220 ;
        RECT 26.700 120.200 26.840 121.920 ;
        RECT 26.640 119.880 26.900 120.200 ;
        RECT 25.260 119.200 25.520 119.520 ;
        RECT 22.500 118.180 22.760 118.500 ;
        RECT 23.420 117.840 23.680 118.160 ;
        RECT 23.480 115.780 23.620 117.840 ;
        RECT 25.320 117.820 25.460 119.200 ;
        RECT 25.260 117.500 25.520 117.820 ;
        RECT 25.720 117.160 25.980 117.480 ;
        RECT 23.420 115.460 23.680 115.780 ;
        RECT 25.780 115.180 25.920 117.160 ;
        RECT 28.480 116.480 28.740 116.800 ;
        RECT 25.780 115.100 26.380 115.180 ;
        RECT 25.720 115.040 26.380 115.100 ;
        RECT 25.720 114.780 25.980 115.040 ;
        RECT 21.120 114.440 21.380 114.760 ;
        RECT 16.800 113.225 18.680 113.595 ;
        RECT 21.120 112.400 21.380 112.720 ;
        RECT 14.220 111.720 14.480 112.040 ;
        RECT 14.280 89.420 14.420 111.720 ;
        RECT 21.180 110.340 21.320 112.400 ;
        RECT 26.240 112.380 26.380 115.040 ;
        RECT 28.540 114.420 28.680 116.480 ;
        RECT 28.480 114.100 28.740 114.420 ;
        RECT 26.180 112.060 26.440 112.380 ;
        RECT 27.560 111.040 27.820 111.360 ;
        RECT 27.620 110.340 27.760 111.040 ;
        RECT 21.120 110.020 21.380 110.340 ;
        RECT 27.560 110.020 27.820 110.340 ;
        RECT 29.460 109.320 29.600 140.960 ;
        RECT 34.920 139.260 35.180 139.580 ;
        RECT 29.860 138.920 30.120 139.240 ;
        RECT 30.320 138.920 30.580 139.240 ;
        RECT 29.920 134.140 30.060 138.920 ;
        RECT 30.380 136.180 30.520 138.920 ;
        RECT 34.460 138.240 34.720 138.560 ;
        RECT 31.800 137.705 33.680 138.075 ;
        RECT 34.520 137.540 34.660 138.240 ;
        RECT 34.460 137.220 34.720 137.540 ;
        RECT 34.000 136.880 34.260 137.200 ;
        RECT 31.240 136.540 31.500 136.860 ;
        RECT 30.320 135.860 30.580 136.180 ;
        RECT 30.780 135.520 31.040 135.840 ;
        RECT 29.860 133.820 30.120 134.140 ;
        RECT 29.920 128.700 30.060 133.820 ;
        RECT 30.840 132.100 30.980 135.520 ;
        RECT 31.300 134.140 31.440 136.540 ;
        RECT 33.540 136.200 33.800 136.520 ;
        RECT 32.620 135.520 32.880 135.840 ;
        RECT 32.680 134.140 32.820 135.520 ;
        RECT 31.240 133.820 31.500 134.140 ;
        RECT 32.160 133.820 32.420 134.140 ;
        RECT 32.620 133.820 32.880 134.140 ;
        RECT 32.220 133.540 32.360 133.820 ;
        RECT 33.600 133.540 33.740 136.200 ;
        RECT 34.060 134.820 34.200 136.880 ;
        RECT 34.980 136.520 35.120 139.260 ;
        RECT 35.440 136.860 35.580 170.880 ;
        RECT 35.900 170.800 36.500 170.940 ;
        RECT 35.900 169.160 36.040 170.800 ;
        RECT 35.840 168.840 36.100 169.160 ;
        RECT 35.900 167.120 36.040 168.840 ;
        RECT 36.820 168.480 36.960 177.000 ;
        RECT 37.280 172.560 37.420 179.720 ;
        RECT 37.740 174.940 37.880 182.780 ;
        RECT 38.200 182.760 38.340 185.500 ;
        RECT 38.140 182.440 38.400 182.760 ;
        RECT 38.200 177.320 38.340 182.440 ;
        RECT 39.520 181.760 39.780 182.080 ;
        RECT 39.580 178.340 39.720 181.760 ;
        RECT 40.900 179.950 41.160 180.040 ;
        RECT 41.420 179.950 41.560 185.500 ;
        RECT 43.660 184.480 43.920 184.800 ;
        RECT 44.120 184.480 44.380 184.800 ;
        RECT 43.720 182.760 43.860 184.480 ;
        RECT 44.180 183.100 44.320 184.480 ;
        RECT 45.100 183.780 45.240 190.600 ;
        RECT 46.020 186.500 46.160 193.660 ;
        RECT 49.180 193.320 49.440 193.640 ;
        RECT 46.420 190.940 46.680 191.260 ;
        RECT 46.480 187.940 46.620 190.940 ;
        RECT 49.240 190.580 49.380 193.320 ;
        RECT 49.180 190.260 49.440 190.580 ;
        RECT 46.800 189.385 48.680 189.755 ;
        RECT 46.880 187.940 47.140 188.200 ;
        RECT 46.480 187.880 47.140 187.940 ;
        RECT 46.480 187.800 47.080 187.880 ;
        RECT 49.240 187.860 49.380 190.260 ;
        RECT 45.960 186.180 46.220 186.500 ;
        RECT 46.480 186.160 46.620 187.800 ;
        RECT 49.180 187.540 49.440 187.860 ;
        RECT 46.420 185.840 46.680 186.160 ;
        RECT 45.500 185.160 45.760 185.480 ;
        RECT 45.040 183.460 45.300 183.780 ;
        RECT 44.120 182.780 44.380 183.100 ;
        RECT 43.660 182.440 43.920 182.760 ;
        RECT 45.560 181.060 45.700 185.160 ;
        RECT 45.960 184.480 46.220 184.800 ;
        RECT 46.420 184.480 46.680 184.800 ;
        RECT 46.020 182.080 46.160 184.480 ;
        RECT 46.480 183.100 46.620 184.480 ;
        RECT 46.800 183.945 48.680 184.315 ;
        RECT 46.420 182.780 46.680 183.100 ;
        RECT 45.960 181.760 46.220 182.080 ;
        RECT 45.500 180.740 45.760 181.060 ;
        RECT 46.480 180.380 46.620 182.780 ;
        RECT 47.340 181.760 47.600 182.080 ;
        RECT 46.880 180.740 47.140 181.060 ;
        RECT 46.940 180.380 47.080 180.740 ;
        RECT 47.400 180.380 47.540 181.760 ;
        RECT 46.420 180.060 46.680 180.380 ;
        RECT 46.880 180.060 47.140 180.380 ;
        RECT 47.340 180.060 47.600 180.380 ;
        RECT 40.430 179.525 40.710 179.895 ;
        RECT 40.900 179.810 41.560 179.950 ;
        RECT 40.900 179.720 41.160 179.810 ;
        RECT 41.810 179.525 42.090 179.895 ;
        RECT 44.120 179.720 44.380 180.040 ;
        RECT 45.500 179.720 45.760 180.040 ;
        RECT 40.500 179.360 40.640 179.525 ;
        RECT 39.980 179.040 40.240 179.360 ;
        RECT 40.440 179.040 40.700 179.360 ;
        RECT 40.900 179.040 41.160 179.360 ;
        RECT 39.520 178.020 39.780 178.340 ;
        RECT 38.140 177.000 38.400 177.320 ;
        RECT 38.200 175.620 38.340 177.000 ;
        RECT 38.140 175.300 38.400 175.620 ;
        RECT 40.040 175.135 40.180 179.040 ;
        RECT 40.960 175.620 41.100 179.040 ;
        RECT 40.900 175.300 41.160 175.620 ;
        RECT 37.680 174.620 37.940 174.940 ;
        RECT 39.970 174.765 40.250 175.135 ;
        RECT 40.440 174.960 40.700 175.280 ;
        RECT 40.040 174.600 40.180 174.765 ;
        RECT 38.140 174.280 38.400 174.600 ;
        RECT 39.980 174.280 40.240 174.600 ;
        RECT 37.220 172.240 37.480 172.560 ;
        RECT 38.200 172.220 38.340 174.280 ;
        RECT 39.060 173.940 39.320 174.260 ;
        RECT 39.520 173.940 39.780 174.260 ;
        RECT 38.140 171.900 38.400 172.220 ;
        RECT 36.760 168.160 37.020 168.480 ;
        RECT 35.840 166.800 36.100 167.120 ;
        RECT 36.820 166.780 36.960 168.160 ;
        RECT 36.760 166.460 37.020 166.780 ;
        RECT 36.820 164.060 36.960 166.460 ;
        RECT 38.140 165.440 38.400 165.760 ;
        RECT 36.760 163.740 37.020 164.060 ;
        RECT 38.200 163.720 38.340 165.440 ;
        RECT 38.140 163.400 38.400 163.720 ;
        RECT 35.840 162.720 36.100 163.040 ;
        RECT 36.300 162.720 36.560 163.040 ;
        RECT 35.900 158.280 36.040 162.720 ;
        RECT 36.360 161.680 36.500 162.720 ;
        RECT 36.300 161.360 36.560 161.680 ;
        RECT 35.840 157.960 36.100 158.280 ;
        RECT 36.360 157.940 36.500 161.360 ;
        RECT 37.680 160.340 37.940 160.660 ;
        RECT 36.300 157.620 36.560 157.940 ;
        RECT 35.840 154.560 36.100 154.880 ;
        RECT 35.900 150.460 36.040 154.560 ;
        RECT 37.740 153.180 37.880 160.340 ;
        RECT 37.220 152.860 37.480 153.180 ;
        RECT 37.680 152.860 37.940 153.180 ;
        RECT 36.760 152.750 37.020 152.840 ;
        RECT 36.360 152.610 37.020 152.750 ;
        RECT 35.840 150.140 36.100 150.460 ;
        RECT 36.360 150.120 36.500 152.610 ;
        RECT 36.760 152.520 37.020 152.610 ;
        RECT 37.280 151.140 37.420 152.860 ;
        RECT 37.220 150.820 37.480 151.140 ;
        RECT 36.300 149.800 36.560 150.120 ;
        RECT 35.840 148.100 36.100 148.420 ;
        RECT 35.900 147.400 36.040 148.100 ;
        RECT 35.840 147.080 36.100 147.400 ;
        RECT 36.360 144.680 36.500 149.800 ;
        RECT 36.760 146.400 37.020 146.720 ;
        RECT 38.600 146.400 38.860 146.720 ;
        RECT 36.300 144.360 36.560 144.680 ;
        RECT 35.840 142.660 36.100 142.980 ;
        RECT 35.900 140.260 36.040 142.660 ;
        RECT 35.840 139.940 36.100 140.260 ;
        RECT 35.840 139.260 36.100 139.580 ;
        RECT 35.380 136.540 35.640 136.860 ;
        RECT 34.920 136.200 35.180 136.520 ;
        RECT 34.460 135.520 34.720 135.840 ;
        RECT 34.000 134.500 34.260 134.820 ;
        RECT 32.220 133.400 34.200 133.540 ;
        RECT 31.240 132.800 31.500 133.120 ;
        RECT 30.780 131.780 31.040 132.100 ;
        RECT 29.860 128.380 30.120 128.700 ;
        RECT 30.320 128.380 30.580 128.700 ;
        RECT 30.380 125.980 30.520 128.380 ;
        RECT 30.320 125.660 30.580 125.980 ;
        RECT 30.780 119.540 31.040 119.860 ;
        RECT 30.840 115.780 30.980 119.540 ;
        RECT 30.780 115.460 31.040 115.780 ;
        RECT 31.300 109.660 31.440 132.800 ;
        RECT 31.800 132.265 33.680 132.635 ;
        RECT 34.060 132.100 34.200 133.400 ;
        RECT 34.000 131.780 34.260 132.100 ;
        RECT 34.000 130.420 34.260 130.740 ;
        RECT 34.060 129.380 34.200 130.420 ;
        RECT 34.000 129.060 34.260 129.380 ;
        RECT 31.800 126.825 33.680 127.195 ;
        RECT 31.800 121.385 33.680 121.755 ;
        RECT 31.800 115.945 33.680 116.315 ;
        RECT 31.800 110.505 33.680 110.875 ;
        RECT 31.240 109.340 31.500 109.660 ;
        RECT 34.520 109.320 34.660 135.520 ;
        RECT 34.920 133.140 35.180 133.460 ;
        RECT 34.980 123.260 35.120 133.140 ;
        RECT 35.900 133.120 36.040 139.260 ;
        RECT 36.360 134.480 36.500 144.360 ;
        RECT 36.820 136.520 36.960 146.400 ;
        RECT 38.140 137.220 38.400 137.540 ;
        RECT 36.760 136.200 37.020 136.520 ;
        RECT 36.300 134.160 36.560 134.480 ;
        RECT 35.840 132.800 36.100 133.120 ;
        RECT 36.360 131.420 36.500 134.160 ;
        RECT 36.300 131.100 36.560 131.420 ;
        RECT 37.680 131.100 37.940 131.420 ;
        RECT 37.740 129.380 37.880 131.100 ;
        RECT 37.680 129.060 37.940 129.380 ;
        RECT 35.840 125.660 36.100 125.980 ;
        RECT 34.920 122.940 35.180 123.260 ;
        RECT 34.980 121.220 35.120 122.940 ;
        RECT 34.920 120.900 35.180 121.220 ;
        RECT 35.900 120.540 36.040 125.660 ;
        RECT 38.200 125.640 38.340 137.220 ;
        RECT 38.660 136.520 38.800 146.400 ;
        RECT 39.120 136.860 39.260 173.940 ;
        RECT 39.580 172.220 39.720 173.940 ;
        RECT 39.520 171.900 39.780 172.220 ;
        RECT 39.980 154.560 40.240 154.880 ;
        RECT 39.520 141.300 39.780 141.620 ;
        RECT 39.580 140.260 39.720 141.300 ;
        RECT 39.520 139.940 39.780 140.260 ;
        RECT 40.040 139.240 40.180 154.560 ;
        RECT 39.980 138.920 40.240 139.240 ;
        RECT 39.060 136.540 39.320 136.860 ;
        RECT 38.600 136.200 38.860 136.520 ;
        RECT 38.600 135.520 38.860 135.840 ;
        RECT 36.760 125.320 37.020 125.640 ;
        RECT 38.140 125.320 38.400 125.640 ;
        RECT 36.820 122.920 36.960 125.320 ;
        RECT 36.760 122.830 37.020 122.920 ;
        RECT 36.360 122.690 37.020 122.830 ;
        RECT 35.840 120.220 36.100 120.540 ;
        RECT 34.920 119.540 35.180 119.860 ;
        RECT 34.980 113.060 35.120 119.540 ;
        RECT 36.360 118.500 36.500 122.690 ;
        RECT 36.760 122.600 37.020 122.690 ;
        RECT 36.760 121.920 37.020 122.240 ;
        RECT 36.300 118.180 36.560 118.500 ;
        RECT 35.380 117.840 35.640 118.160 ;
        RECT 35.440 115.780 35.580 117.840 ;
        RECT 35.380 115.460 35.640 115.780 ;
        RECT 36.820 114.760 36.960 121.920 ;
        RECT 37.680 119.880 37.940 120.200 ;
        RECT 37.740 115.780 37.880 119.880 ;
        RECT 37.680 115.460 37.940 115.780 ;
        RECT 35.840 114.440 36.100 114.760 ;
        RECT 36.760 114.440 37.020 114.760 ;
        RECT 35.900 114.080 36.040 114.440 ;
        RECT 35.840 113.760 36.100 114.080 ;
        RECT 34.920 112.740 35.180 113.060 ;
        RECT 35.900 112.380 36.040 113.760 ;
        RECT 35.840 112.060 36.100 112.380 ;
        RECT 36.760 111.380 37.020 111.700 ;
        RECT 29.400 109.000 29.660 109.320 ;
        RECT 34.460 109.000 34.720 109.320 ;
        RECT 27.560 108.660 27.820 108.980 ;
        RECT 23.420 108.320 23.680 108.640 ;
        RECT 16.800 107.785 18.680 108.155 ;
        RECT 23.480 107.280 23.620 108.320 ;
        RECT 23.420 106.960 23.680 107.280 ;
        RECT 18.820 106.280 19.080 106.600 ;
        RECT 16.800 102.345 18.680 102.715 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 18.880 88.660 19.020 106.280 ;
        RECT 27.620 103.880 27.760 108.660 ;
        RECT 31.700 108.320 31.960 108.640 ;
        RECT 32.160 108.320 32.420 108.640 ;
        RECT 34.000 108.320 34.260 108.640 ;
        RECT 31.760 107.280 31.900 108.320 ;
        RECT 32.220 107.620 32.360 108.320 ;
        RECT 32.160 107.300 32.420 107.620 ;
        RECT 31.700 106.960 31.960 107.280 ;
        RECT 28.940 106.280 29.200 106.600 ;
        RECT 30.320 106.280 30.580 106.600 ;
        RECT 29.000 104.900 29.140 106.280 ;
        RECT 28.940 104.580 29.200 104.900 ;
        RECT 27.560 103.560 27.820 103.880 ;
        RECT 28.020 102.880 28.280 103.200 ;
        RECT 28.080 101.500 28.220 102.880 ;
        RECT 28.020 101.180 28.280 101.500 ;
        RECT 26.180 100.840 26.440 101.160 ;
        RECT 19.910 88.660 21.130 89.850 ;
        RECT 26.240 89.210 26.380 100.840 ;
        RECT 26.170 88.990 26.450 89.210 ;
        RECT 18.880 88.520 21.130 88.660 ;
        RECT 19.910 85.980 21.130 88.520 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 30.380 88.660 30.520 106.280 ;
        RECT 31.800 105.065 33.680 105.435 ;
        RECT 34.060 101.840 34.200 108.320 ;
        RECT 36.820 106.940 36.960 111.380 ;
        RECT 38.660 106.940 38.800 135.520 ;
        RECT 40.500 134.140 40.640 174.960 ;
        RECT 40.960 172.220 41.100 175.300 ;
        RECT 41.880 174.260 42.020 179.525 ;
        RECT 42.280 179.040 42.540 179.360 ;
        RECT 41.820 173.940 42.080 174.260 ;
        RECT 40.900 171.900 41.160 172.220 ;
        RECT 40.960 169.840 41.100 171.900 ;
        RECT 41.360 170.880 41.620 171.200 ;
        RECT 40.900 169.520 41.160 169.840 ;
        RECT 40.960 156.240 41.100 169.520 ;
        RECT 40.900 155.920 41.160 156.240 ;
        RECT 40.900 149.120 41.160 149.440 ;
        RECT 40.960 134.140 41.100 149.120 ;
        RECT 41.420 139.920 41.560 170.880 ;
        RECT 42.340 160.180 42.480 179.040 ;
        RECT 43.660 177.340 43.920 177.660 ;
        RECT 42.740 176.320 43.000 176.640 ;
        RECT 42.800 172.220 42.940 176.320 ;
        RECT 43.720 174.600 43.860 177.340 ;
        RECT 44.180 174.600 44.320 179.720 ;
        RECT 44.580 179.040 44.840 179.360 ;
        RECT 44.640 174.600 44.780 179.040 ;
        RECT 45.560 177.660 45.700 179.720 ;
        RECT 46.940 179.610 47.080 180.060 ;
        RECT 46.480 179.470 47.080 179.610 ;
        RECT 45.960 179.040 46.220 179.360 ;
        RECT 46.020 178.340 46.160 179.040 ;
        RECT 45.960 178.020 46.220 178.340 ;
        RECT 45.500 177.340 45.760 177.660 ;
        RECT 45.560 174.940 45.700 177.340 ;
        RECT 46.480 175.620 46.620 179.470 ;
        RECT 46.800 178.505 48.680 178.875 ;
        RECT 47.800 177.340 48.060 177.660 ;
        RECT 49.180 177.340 49.440 177.660 ;
        RECT 46.420 175.300 46.680 175.620 ;
        RECT 45.500 174.620 45.760 174.940 ;
        RECT 43.660 174.280 43.920 174.600 ;
        RECT 44.120 174.280 44.380 174.600 ;
        RECT 44.580 174.280 44.840 174.600 ;
        RECT 44.640 172.900 44.780 174.280 ;
        RECT 47.860 174.260 48.000 177.340 ;
        RECT 45.500 173.940 45.760 174.260 ;
        RECT 47.800 173.940 48.060 174.260 ;
        RECT 44.580 172.580 44.840 172.900 ;
        RECT 42.740 171.900 43.000 172.220 ;
        RECT 44.110 169.325 44.390 169.695 ;
        RECT 44.180 169.160 44.320 169.325 ;
        RECT 44.120 168.840 44.380 169.160 ;
        RECT 43.200 166.120 43.460 166.440 ;
        RECT 42.740 165.440 43.000 165.760 ;
        RECT 42.800 162.020 42.940 165.440 ;
        RECT 42.740 161.700 43.000 162.020 ;
        RECT 42.340 160.040 42.940 160.180 ;
        RECT 41.820 157.960 42.080 158.280 ;
        RECT 41.880 156.580 42.020 157.960 ;
        RECT 42.280 157.280 42.540 157.600 ;
        RECT 41.820 156.260 42.080 156.580 ;
        RECT 41.810 155.725 42.090 156.095 ;
        RECT 41.820 155.580 42.080 155.725 ;
        RECT 41.820 151.840 42.080 152.160 ;
        RECT 41.880 150.460 42.020 151.840 ;
        RECT 41.820 150.140 42.080 150.460 ;
        RECT 41.880 146.720 42.020 150.140 ;
        RECT 41.820 146.400 42.080 146.720 ;
        RECT 41.360 139.600 41.620 139.920 ;
        RECT 42.340 136.520 42.480 157.280 ;
        RECT 42.280 136.200 42.540 136.520 ;
        RECT 42.800 134.140 42.940 160.040 ;
        RECT 43.260 158.280 43.400 166.120 ;
        RECT 43.200 157.960 43.460 158.280 ;
        RECT 45.040 157.960 45.300 158.280 ;
        RECT 43.200 157.280 43.460 157.600 ;
        RECT 43.260 156.095 43.400 157.280 ;
        RECT 45.100 156.580 45.240 157.960 ;
        RECT 45.040 156.260 45.300 156.580 ;
        RECT 43.190 155.725 43.470 156.095 ;
        RECT 43.260 155.470 43.400 155.725 ;
        RECT 43.660 155.470 43.920 155.560 ;
        RECT 43.260 155.330 43.920 155.470 ;
        RECT 43.660 155.240 43.920 155.330 ;
        RECT 43.660 154.560 43.920 154.880 ;
        RECT 45.040 154.560 45.300 154.880 ;
        RECT 43.200 152.180 43.460 152.500 ;
        RECT 43.260 150.460 43.400 152.180 ;
        RECT 43.200 150.140 43.460 150.460 ;
        RECT 43.260 147.060 43.400 150.140 ;
        RECT 43.200 146.740 43.460 147.060 ;
        RECT 43.720 134.140 43.860 154.560 ;
        RECT 44.580 152.695 44.840 152.840 ;
        RECT 44.570 152.325 44.850 152.695 ;
        RECT 44.120 149.120 44.380 149.440 ;
        RECT 40.440 133.820 40.700 134.140 ;
        RECT 40.900 133.820 41.160 134.140 ;
        RECT 42.740 133.820 43.000 134.140 ;
        RECT 43.660 133.820 43.920 134.140 ;
        RECT 44.180 133.540 44.320 149.120 ;
        RECT 44.640 147.400 44.780 152.325 ;
        RECT 45.100 150.460 45.240 154.560 ;
        RECT 45.040 150.140 45.300 150.460 ;
        RECT 44.580 147.080 44.840 147.400 ;
        RECT 45.040 142.320 45.300 142.640 ;
        RECT 44.580 137.220 44.840 137.540 ;
        RECT 43.720 133.400 44.320 133.540 ;
        RECT 39.520 132.800 39.780 133.120 ;
        RECT 40.440 132.800 40.700 133.120 ;
        RECT 41.360 132.800 41.620 133.120 ;
        RECT 43.200 132.800 43.460 133.120 ;
        RECT 39.580 128.700 39.720 132.800 ;
        RECT 39.980 131.440 40.240 131.760 ;
        RECT 39.520 128.380 39.780 128.700 ;
        RECT 40.040 125.300 40.180 131.440 ;
        RECT 40.500 125.640 40.640 132.800 ;
        RECT 40.440 125.320 40.700 125.640 ;
        RECT 39.980 124.980 40.240 125.300 ;
        RECT 39.980 119.200 40.240 119.520 ;
        RECT 39.060 117.160 39.320 117.480 ;
        RECT 39.120 115.780 39.260 117.160 ;
        RECT 39.060 115.460 39.320 115.780 ;
        RECT 40.040 114.760 40.180 119.200 ;
        RECT 39.980 114.440 40.240 114.760 ;
        RECT 40.900 108.660 41.160 108.980 ;
        RECT 40.960 107.280 41.100 108.660 ;
        RECT 40.900 106.960 41.160 107.280 ;
        RECT 41.420 106.940 41.560 132.800 ;
        RECT 42.740 130.080 43.000 130.400 ;
        RECT 42.800 129.040 42.940 130.080 ;
        RECT 42.740 128.720 43.000 129.040 ;
        RECT 42.740 128.040 43.000 128.360 ;
        RECT 42.280 125.320 42.540 125.640 ;
        RECT 41.820 122.600 42.080 122.920 ;
        RECT 41.880 120.200 42.020 122.600 ;
        RECT 41.820 119.880 42.080 120.200 ;
        RECT 42.340 119.520 42.480 125.320 ;
        RECT 42.800 123.940 42.940 128.040 ;
        RECT 43.260 125.300 43.400 132.800 ;
        RECT 43.720 129.380 43.860 133.400 ;
        RECT 44.120 132.800 44.380 133.120 ;
        RECT 43.660 129.060 43.920 129.380 ;
        RECT 43.200 124.980 43.460 125.300 ;
        RECT 42.740 123.620 43.000 123.940 ;
        RECT 43.660 122.260 43.920 122.580 ;
        RECT 43.720 120.540 43.860 122.260 ;
        RECT 43.660 120.220 43.920 120.540 ;
        RECT 42.280 119.200 42.540 119.520 ;
        RECT 42.340 118.500 42.480 119.200 ;
        RECT 42.280 118.180 42.540 118.500 ;
        RECT 42.340 114.420 42.480 118.180 ;
        RECT 43.200 117.840 43.460 118.160 ;
        RECT 43.260 115.780 43.400 117.840 ;
        RECT 43.200 115.460 43.460 115.780 ;
        RECT 43.720 115.440 43.860 120.220 ;
        RECT 43.660 115.120 43.920 115.440 ;
        RECT 42.280 114.100 42.540 114.420 ;
        RECT 44.180 111.880 44.320 132.800 ;
        RECT 44.640 125.640 44.780 137.220 ;
        RECT 45.100 129.380 45.240 142.320 ;
        RECT 45.560 136.860 45.700 173.940 ;
        RECT 46.800 173.065 48.680 173.435 ;
        RECT 49.240 172.900 49.380 177.340 ;
        RECT 49.700 172.900 49.840 194.430 ;
        RECT 50.560 194.340 50.820 194.430 ;
        RECT 53.380 194.320 53.520 195.360 ;
        RECT 53.320 194.000 53.580 194.320 ;
        RECT 50.560 193.320 50.820 193.640 ;
        RECT 50.620 191.940 50.760 193.320 ;
        RECT 54.240 192.640 54.500 192.960 ;
        RECT 50.560 191.620 50.820 191.940 ;
        RECT 52.400 190.940 52.660 191.260 ;
        RECT 50.100 187.200 50.360 187.520 ;
        RECT 50.160 183.780 50.300 187.200 ;
        RECT 50.100 183.460 50.360 183.780 ;
        RECT 50.100 182.440 50.360 182.760 ;
        RECT 50.160 181.060 50.300 182.440 ;
        RECT 50.100 180.740 50.360 181.060 ;
        RECT 52.460 180.380 52.600 190.940 ;
        RECT 54.300 190.920 54.440 192.640 ;
        RECT 54.240 190.600 54.500 190.920 ;
        RECT 57.980 190.240 58.120 195.360 ;
        RECT 61.800 192.105 63.680 192.475 ;
        RECT 63.960 191.600 64.100 202.500 ;
        RECT 64.880 201.460 65.020 203.520 ;
        RECT 64.820 201.140 65.080 201.460 ;
        RECT 64.820 198.080 65.080 198.400 ;
        RECT 63.900 191.280 64.160 191.600 ;
        RECT 59.300 190.940 59.560 191.260 ;
        RECT 57.920 189.920 58.180 190.240 ;
        RECT 57.980 189.220 58.120 189.920 ;
        RECT 57.920 188.900 58.180 189.220 ;
        RECT 55.620 188.220 55.880 188.540 ;
        RECT 56.540 188.220 56.800 188.540 ;
        RECT 55.680 188.055 55.820 188.220 ;
        RECT 55.610 187.685 55.890 188.055 ;
        RECT 56.080 181.760 56.340 182.080 ;
        RECT 52.400 180.060 52.660 180.380 ;
        RECT 54.240 180.060 54.500 180.380 ;
        RECT 50.560 179.040 50.820 179.360 ;
        RECT 50.620 177.660 50.760 179.040 ;
        RECT 52.460 178.000 52.600 180.060 ;
        RECT 53.780 179.380 54.040 179.700 ;
        RECT 53.840 178.340 53.980 179.380 ;
        RECT 53.780 178.020 54.040 178.340 ;
        RECT 52.400 177.680 52.660 178.000 ;
        RECT 50.560 177.340 50.820 177.660 ;
        RECT 51.020 176.660 51.280 176.980 ;
        RECT 50.100 176.320 50.360 176.640 ;
        RECT 49.180 172.580 49.440 172.900 ;
        RECT 49.640 172.580 49.900 172.900 ;
        RECT 49.240 172.220 49.380 172.580 ;
        RECT 47.340 171.900 47.600 172.220 ;
        RECT 49.180 171.900 49.440 172.220 ;
        RECT 49.640 171.900 49.900 172.220 ;
        RECT 45.960 170.880 46.220 171.200 ;
        RECT 46.020 160.180 46.160 170.880 ;
        RECT 47.400 170.180 47.540 171.900 ;
        RECT 49.700 171.540 49.840 171.900 ;
        RECT 49.640 171.220 49.900 171.540 ;
        RECT 47.340 169.860 47.600 170.180 ;
        RECT 46.800 167.625 48.680 167.995 ;
        RECT 49.640 165.440 49.900 165.760 ;
        RECT 49.180 163.400 49.440 163.720 ;
        RECT 46.420 163.060 46.680 163.380 ;
        RECT 46.480 162.020 46.620 163.060 ;
        RECT 46.800 162.185 48.680 162.555 ;
        RECT 49.240 162.020 49.380 163.400 ;
        RECT 49.700 162.020 49.840 165.440 ;
        RECT 46.420 161.700 46.680 162.020 ;
        RECT 49.180 161.700 49.440 162.020 ;
        RECT 49.640 161.700 49.900 162.020 ;
        RECT 49.640 161.020 49.900 161.340 ;
        RECT 49.180 160.680 49.440 161.000 ;
        RECT 46.020 160.040 46.620 160.180 ;
        RECT 45.960 157.280 46.220 157.600 ;
        RECT 46.020 141.960 46.160 157.280 ;
        RECT 46.480 142.300 46.620 160.040 ;
        RECT 46.800 156.745 48.680 157.115 ;
        RECT 49.240 156.580 49.380 160.680 ;
        RECT 49.700 159.300 49.840 161.020 ;
        RECT 49.640 158.980 49.900 159.300 ;
        RECT 50.160 158.020 50.300 176.320 ;
        RECT 51.080 172.900 51.220 176.660 ;
        RECT 54.300 175.620 54.440 180.060 ;
        RECT 56.140 178.000 56.280 181.760 ;
        RECT 56.600 180.720 56.740 188.220 ;
        RECT 59.360 187.860 59.500 190.940 ;
        RECT 60.220 190.260 60.480 190.580 ;
        RECT 60.280 189.220 60.420 190.260 ;
        RECT 62.060 189.920 62.320 190.240 ;
        RECT 60.220 188.900 60.480 189.220 ;
        RECT 62.120 188.200 62.260 189.920 ;
        RECT 62.060 187.880 62.320 188.200 ;
        RECT 59.300 187.540 59.560 187.860 ;
        RECT 59.360 185.820 59.500 187.540 ;
        RECT 64.880 187.260 65.020 198.080 ;
        RECT 66.260 193.980 66.400 204.540 ;
        RECT 73.160 203.840 73.300 206.920 ;
        RECT 73.100 203.520 73.360 203.840 ;
        RECT 66.660 202.500 66.920 202.820 ;
        RECT 66.200 193.660 66.460 193.980 ;
        RECT 65.740 192.640 66.000 192.960 ;
        RECT 65.800 190.580 65.940 192.640 ;
        RECT 65.740 190.260 66.000 190.580 ;
        RECT 66.260 190.240 66.400 193.660 ;
        RECT 66.200 189.920 66.460 190.240 ;
        RECT 65.740 187.880 66.000 188.200 ;
        RECT 64.420 187.120 65.020 187.260 ;
        RECT 61.800 186.665 63.680 187.035 ;
        RECT 60.680 185.840 60.940 186.160 ;
        RECT 59.300 185.500 59.560 185.820 ;
        RECT 57.920 184.820 58.180 185.140 ;
        RECT 57.980 183.780 58.120 184.820 ;
        RECT 57.920 183.460 58.180 183.780 ;
        RECT 59.360 183.100 59.500 185.500 ;
        RECT 60.740 183.100 60.880 185.840 ;
        RECT 59.300 182.780 59.560 183.100 ;
        RECT 60.680 182.780 60.940 183.100 ;
        RECT 56.540 180.400 56.800 180.720 ;
        RECT 56.080 177.680 56.340 178.000 ;
        RECT 54.240 175.300 54.500 175.620 ;
        RECT 54.300 174.940 54.440 175.300 ;
        RECT 53.780 174.620 54.040 174.940 ;
        RECT 54.240 174.620 54.500 174.940 ;
        RECT 53.320 173.940 53.580 174.260 ;
        RECT 51.020 172.580 51.280 172.900 ;
        RECT 51.080 172.220 51.220 172.580 ;
        RECT 53.380 172.220 53.520 173.940 ;
        RECT 53.840 172.220 53.980 174.620 ;
        RECT 56.600 174.600 56.740 180.400 ;
        RECT 57.920 179.040 58.180 179.360 ;
        RECT 57.980 174.940 58.120 179.040 ;
        RECT 59.360 177.320 59.500 182.780 ;
        RECT 59.300 177.000 59.560 177.320 ;
        RECT 57.920 174.620 58.180 174.940 ;
        RECT 54.690 174.085 54.970 174.455 ;
        RECT 56.540 174.280 56.800 174.600 ;
        RECT 54.760 172.900 54.900 174.085 ;
        RECT 57.000 173.600 57.260 173.920 ;
        RECT 54.700 172.580 54.960 172.900 ;
        RECT 54.760 172.220 54.900 172.580 ;
        RECT 57.060 172.560 57.200 173.600 ;
        RECT 57.000 172.240 57.260 172.560 ;
        RECT 60.740 172.220 60.880 182.780 ;
        RECT 61.800 181.225 63.680 181.595 ;
        RECT 61.200 178.340 62.260 178.420 ;
        RECT 61.200 178.280 62.320 178.340 ;
        RECT 61.200 178.000 61.340 178.280 ;
        RECT 62.060 178.020 62.320 178.280 ;
        RECT 61.140 177.680 61.400 178.000 ;
        RECT 63.900 177.000 64.160 177.320 ;
        RECT 61.800 175.785 63.680 176.155 ;
        RECT 63.960 175.620 64.100 177.000 ;
        RECT 63.900 175.300 64.160 175.620 ;
        RECT 61.140 173.940 61.400 174.260 ;
        RECT 62.970 174.085 63.250 174.455 ;
        RECT 61.200 172.900 61.340 173.940 ;
        RECT 63.040 173.920 63.180 174.085 ;
        RECT 62.980 173.600 63.240 173.920 ;
        RECT 61.140 172.580 61.400 172.900 ;
        RECT 51.020 171.900 51.280 172.220 ;
        RECT 53.320 171.900 53.580 172.220 ;
        RECT 53.780 171.900 54.040 172.220 ;
        RECT 54.700 171.900 54.960 172.220 ;
        RECT 60.680 171.900 60.940 172.220 ;
        RECT 52.400 170.880 52.660 171.200 ;
        RECT 51.020 166.800 51.280 167.120 ;
        RECT 51.080 164.740 51.220 166.800 ;
        RECT 51.020 164.420 51.280 164.740 ;
        RECT 50.560 158.980 50.820 159.300 ;
        RECT 50.620 158.620 50.760 158.980 ;
        RECT 50.560 158.300 50.820 158.620 ;
        RECT 49.700 157.880 50.300 158.020 ;
        RECT 49.180 156.260 49.440 156.580 ;
        RECT 46.880 155.580 47.140 155.900 ;
        RECT 46.940 155.220 47.080 155.580 ;
        RECT 46.880 154.900 47.140 155.220 ;
        RECT 49.180 154.560 49.440 154.880 ;
        RECT 46.800 151.305 48.680 151.675 ;
        RECT 49.240 150.540 49.380 154.560 ;
        RECT 48.780 150.400 49.380 150.540 ;
        RECT 49.700 150.460 49.840 157.880 ;
        RECT 50.100 157.280 50.360 157.600 ;
        RECT 50.160 150.460 50.300 157.280 ;
        RECT 50.560 156.260 50.820 156.580 ;
        RECT 50.620 152.160 50.760 156.260 ;
        RECT 51.020 152.520 51.280 152.840 ;
        RECT 50.560 151.840 50.820 152.160 ;
        RECT 48.780 147.400 48.920 150.400 ;
        RECT 49.640 150.140 49.900 150.460 ;
        RECT 50.100 150.140 50.360 150.460 ;
        RECT 50.560 149.800 50.820 150.120 ;
        RECT 50.620 148.420 50.760 149.800 ;
        RECT 49.180 148.100 49.440 148.420 ;
        RECT 50.560 148.100 50.820 148.420 ;
        RECT 48.720 147.080 48.980 147.400 ;
        RECT 46.800 145.865 48.680 146.235 ;
        RECT 49.240 144.420 49.380 148.100 ;
        RECT 49.640 146.400 49.900 146.720 ;
        RECT 49.700 145.020 49.840 146.400 ;
        RECT 51.080 145.700 51.220 152.520 ;
        RECT 51.480 149.120 51.740 149.440 ;
        RECT 51.540 147.060 51.680 149.120 ;
        RECT 52.460 147.740 52.600 170.880 ;
        RECT 53.320 166.800 53.580 167.120 ;
        RECT 53.380 163.720 53.520 166.800 ;
        RECT 54.240 166.120 54.500 166.440 ;
        RECT 54.700 166.120 54.960 166.440 ;
        RECT 57.460 166.120 57.720 166.440 ;
        RECT 53.320 163.400 53.580 163.720 ;
        RECT 52.860 162.720 53.120 163.040 ;
        RECT 52.920 159.300 53.060 162.720 ;
        RECT 54.300 162.020 54.440 166.120 ;
        RECT 54.760 164.740 54.900 166.120 ;
        RECT 54.700 164.420 54.960 164.740 ;
        RECT 57.520 164.400 57.660 166.120 ;
        RECT 58.840 165.440 59.100 165.760 ;
        RECT 57.460 164.080 57.720 164.400 ;
        RECT 58.900 163.380 59.040 165.440 ;
        RECT 60.740 164.060 60.880 171.900 ;
        RECT 61.800 170.345 63.680 170.715 ;
        RECT 61.600 166.460 61.860 166.780 ;
        RECT 61.660 166.180 61.800 166.460 ;
        RECT 61.200 166.040 61.800 166.180 ;
        RECT 63.900 166.120 64.160 166.440 ;
        RECT 61.200 164.140 61.340 166.040 ;
        RECT 61.800 164.905 63.680 165.275 ;
        RECT 61.600 164.420 61.860 164.740 ;
        RECT 61.660 164.140 61.800 164.420 ;
        RECT 60.680 163.740 60.940 164.060 ;
        RECT 61.200 164.000 61.800 164.140 ;
        RECT 58.840 163.060 59.100 163.380 ;
        RECT 54.240 161.700 54.500 162.020 ;
        RECT 53.320 160.340 53.580 160.660 ;
        RECT 52.860 158.980 53.120 159.300 ;
        RECT 52.920 158.280 53.060 158.980 ;
        RECT 52.860 157.960 53.120 158.280 ;
        RECT 53.380 157.600 53.520 160.340 ;
        RECT 53.780 157.960 54.040 158.280 ;
        RECT 57.000 157.960 57.260 158.280 ;
        RECT 61.200 158.190 61.340 164.000 ;
        RECT 63.960 163.720 64.100 166.120 ;
        RECT 63.900 163.400 64.160 163.720 ;
        RECT 62.520 163.060 62.780 163.380 ;
        RECT 62.580 162.020 62.720 163.060 ;
        RECT 62.520 161.700 62.780 162.020 ;
        RECT 61.800 159.465 63.680 159.835 ;
        RECT 62.980 158.190 63.240 158.280 ;
        RECT 61.200 158.050 63.240 158.190 ;
        RECT 62.980 157.960 63.240 158.050 ;
        RECT 53.320 157.280 53.580 157.600 ;
        RECT 53.380 156.240 53.520 157.280 ;
        RECT 53.320 155.920 53.580 156.240 ;
        RECT 53.840 155.900 53.980 157.960 ;
        RECT 53.780 155.580 54.040 155.900 ;
        RECT 53.780 154.560 54.040 154.880 ;
        RECT 54.240 154.560 54.500 154.880 ;
        RECT 53.840 150.460 53.980 154.560 ;
        RECT 54.300 153.520 54.440 154.560 ;
        RECT 54.240 153.200 54.500 153.520 ;
        RECT 57.060 152.840 57.200 157.960 ;
        RECT 58.840 157.280 59.100 157.600 ;
        RECT 58.900 156.240 59.040 157.280 ;
        RECT 58.840 155.920 59.100 156.240 ;
        RECT 63.960 155.900 64.100 163.400 ;
        RECT 63.900 155.580 64.160 155.900 ;
        RECT 61.140 155.240 61.400 155.560 ;
        RECT 57.000 152.520 57.260 152.840 ;
        RECT 58.840 151.840 59.100 152.160 ;
        RECT 58.900 150.460 59.040 151.840 ;
        RECT 61.200 151.140 61.340 155.240 ;
        RECT 61.800 154.025 63.680 154.395 ;
        RECT 64.420 153.180 64.560 187.120 ;
        RECT 65.800 180.040 65.940 187.880 ;
        RECT 65.740 179.720 66.000 180.040 ;
        RECT 66.200 179.040 66.460 179.360 ;
        RECT 66.260 177.855 66.400 179.040 ;
        RECT 66.190 177.485 66.470 177.855 ;
        RECT 65.280 176.660 65.540 176.980 ;
        RECT 64.820 176.320 65.080 176.640 ;
        RECT 64.880 174.940 65.020 176.320 ;
        RECT 65.340 175.135 65.480 176.660 ;
        RECT 66.200 175.300 66.460 175.620 ;
        RECT 64.820 174.620 65.080 174.940 ;
        RECT 65.270 174.765 65.550 175.135 ;
        RECT 66.260 174.940 66.400 175.300 ;
        RECT 66.200 174.620 66.460 174.940 ;
        RECT 64.820 173.940 65.080 174.260 ;
        RECT 64.880 172.900 65.020 173.940 ;
        RECT 64.820 172.580 65.080 172.900 ;
        RECT 66.720 166.440 66.860 202.500 ;
        RECT 73.160 202.140 73.300 203.520 ;
        RECT 73.100 201.820 73.360 202.140 ;
        RECT 71.720 200.800 71.980 201.120 ;
        RECT 72.640 200.800 72.900 201.120 ;
        RECT 71.780 199.420 71.920 200.800 ;
        RECT 68.500 199.100 68.760 199.420 ;
        RECT 71.720 199.100 71.980 199.420 ;
        RECT 68.560 197.380 68.700 199.100 ;
        RECT 72.700 198.400 72.840 200.800 ;
        RECT 73.620 198.740 73.760 207.600 ;
        RECT 79.540 207.260 79.800 207.580 ;
        RECT 74.020 206.240 74.280 206.560 ;
        RECT 75.860 206.240 76.120 206.560 ;
        RECT 74.080 205.540 74.220 206.240 ;
        RECT 74.020 205.220 74.280 205.540 ;
        RECT 75.920 205.200 76.060 206.240 ;
        RECT 76.800 205.705 78.680 206.075 ;
        RECT 75.860 204.880 76.120 205.200 ;
        RECT 74.020 203.520 74.280 203.840 ;
        RECT 74.080 201.800 74.220 203.520 ;
        RECT 76.320 202.160 76.580 202.480 ;
        RECT 74.480 201.820 74.740 202.140 ;
        RECT 74.020 201.480 74.280 201.800 ;
        RECT 74.080 200.100 74.220 201.480 ;
        RECT 74.020 199.780 74.280 200.100 ;
        RECT 74.540 199.760 74.680 201.820 ;
        RECT 74.940 201.140 75.200 201.460 ;
        RECT 75.400 201.140 75.660 201.460 ;
        RECT 75.000 200.100 75.140 201.140 ;
        RECT 74.940 199.780 75.200 200.100 ;
        RECT 74.480 199.440 74.740 199.760 ;
        RECT 73.100 198.420 73.360 198.740 ;
        RECT 73.560 198.420 73.820 198.740 ;
        RECT 72.640 198.080 72.900 198.400 ;
        RECT 68.500 197.060 68.760 197.380 ;
        RECT 69.880 197.060 70.140 197.380 ;
        RECT 68.960 196.040 69.220 196.360 ;
        RECT 69.020 193.980 69.160 196.040 ;
        RECT 68.960 193.660 69.220 193.980 ;
        RECT 69.940 190.660 70.080 197.060 ;
        RECT 72.700 196.700 72.840 198.080 ;
        RECT 73.160 196.700 73.300 198.420 ;
        RECT 73.620 197.380 73.760 198.420 ;
        RECT 73.560 197.060 73.820 197.380 ;
        RECT 70.340 196.380 70.600 196.700 ;
        RECT 72.640 196.380 72.900 196.700 ;
        RECT 73.100 196.380 73.360 196.700 ;
        RECT 70.400 192.960 70.540 196.380 ;
        RECT 71.720 195.700 71.980 196.020 ;
        RECT 71.780 194.660 71.920 195.700 ;
        RECT 71.720 194.340 71.980 194.660 ;
        RECT 72.700 194.320 72.840 196.380 ;
        RECT 72.640 194.000 72.900 194.320 ;
        RECT 73.160 193.980 73.300 196.380 ;
        RECT 73.100 193.660 73.360 193.980 ;
        RECT 70.340 192.640 70.600 192.960 ;
        RECT 72.640 192.870 72.900 192.960 ;
        RECT 72.240 192.730 72.900 192.870 ;
        RECT 71.260 190.940 71.520 191.260 ;
        RECT 71.320 190.660 71.460 190.940 ;
        RECT 69.940 190.520 71.460 190.660 ;
        RECT 69.880 189.920 70.140 190.240 ;
        RECT 68.040 185.500 68.300 185.820 ;
        RECT 68.100 183.100 68.240 185.500 ;
        RECT 68.040 182.780 68.300 183.100 ;
        RECT 69.420 181.760 69.680 182.080 ;
        RECT 67.580 180.400 67.840 180.720 ;
        RECT 67.640 179.895 67.780 180.400 ;
        RECT 67.570 179.525 67.850 179.895 ;
        RECT 68.500 179.780 68.760 180.040 ;
        RECT 68.500 179.720 69.160 179.780 ;
        RECT 68.560 179.640 69.160 179.720 ;
        RECT 69.020 177.660 69.160 179.640 ;
        RECT 69.480 177.660 69.620 181.760 ;
        RECT 68.960 177.340 69.220 177.660 ;
        RECT 69.420 177.340 69.680 177.660 ;
        RECT 69.020 176.640 69.160 177.340 ;
        RECT 68.040 176.320 68.300 176.640 ;
        RECT 68.960 176.320 69.220 176.640 ;
        RECT 68.100 175.620 68.240 176.320 ;
        RECT 68.040 175.300 68.300 175.620 ;
        RECT 69.940 174.940 70.080 189.920 ;
        RECT 72.240 188.200 72.380 192.730 ;
        RECT 72.640 192.640 72.900 192.730 ;
        RECT 73.160 191.340 73.300 193.660 ;
        RECT 72.700 191.200 73.300 191.340 ;
        RECT 72.180 187.880 72.440 188.200 ;
        RECT 71.260 185.840 71.520 186.160 ;
        RECT 71.320 183.780 71.460 185.840 ;
        RECT 71.260 183.460 71.520 183.780 ;
        RECT 71.720 183.460 71.980 183.780 ;
        RECT 71.780 183.100 71.920 183.460 ;
        RECT 71.720 182.780 71.980 183.100 ;
        RECT 72.240 183.010 72.380 187.880 ;
        RECT 72.700 185.140 72.840 191.200 ;
        RECT 73.100 190.600 73.360 190.920 ;
        RECT 73.160 189.220 73.300 190.600 ;
        RECT 73.620 190.580 73.760 197.060 ;
        RECT 74.540 196.360 74.680 199.440 ;
        RECT 74.480 196.040 74.740 196.360 ;
        RECT 74.540 190.920 74.680 196.040 ;
        RECT 75.460 196.020 75.600 201.140 ;
        RECT 75.860 200.800 76.120 201.120 ;
        RECT 75.920 199.080 76.060 200.800 ;
        RECT 76.380 200.100 76.520 202.160 ;
        RECT 79.080 201.820 79.340 202.140 ;
        RECT 76.800 200.265 78.680 200.635 ;
        RECT 76.320 199.780 76.580 200.100 ;
        RECT 79.140 199.420 79.280 201.820 ;
        RECT 79.600 201.460 79.740 207.260 ;
        RECT 106.800 205.705 108.680 206.075 ;
        RECT 83.680 204.880 83.940 205.200 ;
        RECT 79.540 201.140 79.800 201.460 ;
        RECT 79.600 200.100 79.740 201.140 ;
        RECT 83.740 200.100 83.880 204.880 ;
        RECT 88.280 204.200 88.540 204.520 ;
        RECT 84.600 201.820 84.860 202.140 ;
        RECT 84.660 200.100 84.800 201.820 ;
        RECT 88.340 201.800 88.480 204.200 ;
        RECT 91.800 202.985 93.680 203.355 ;
        RECT 121.800 202.985 123.680 203.355 ;
        RECT 88.280 201.480 88.540 201.800 ;
        RECT 96.560 201.480 96.820 201.800 ;
        RECT 85.520 201.140 85.780 201.460 ;
        RECT 85.580 200.100 85.720 201.140 ;
        RECT 79.540 199.780 79.800 200.100 ;
        RECT 83.680 199.780 83.940 200.100 ;
        RECT 84.600 199.780 84.860 200.100 ;
        RECT 85.520 199.780 85.780 200.100 ;
        RECT 80.920 199.440 81.180 199.760 ;
        RECT 79.080 199.100 79.340 199.420 ;
        RECT 80.000 199.100 80.260 199.420 ;
        RECT 75.860 198.760 76.120 199.080 ;
        RECT 80.060 197.040 80.200 199.100 ;
        RECT 80.980 198.400 81.120 199.440 ;
        RECT 86.900 199.100 87.160 199.420 ;
        RECT 80.920 198.080 81.180 198.400 ;
        RECT 80.000 196.720 80.260 197.040 ;
        RECT 75.400 195.700 75.660 196.020 ;
        RECT 76.800 194.825 78.680 195.195 ;
        RECT 76.320 193.660 76.580 193.980 ;
        RECT 74.480 190.600 74.740 190.920 ;
        RECT 73.560 190.260 73.820 190.580 ;
        RECT 73.100 188.900 73.360 189.220 ;
        RECT 73.620 185.820 73.760 190.260 ;
        RECT 73.560 185.500 73.820 185.820 ;
        RECT 72.640 184.820 72.900 185.140 ;
        RECT 72.700 183.780 72.840 184.820 ;
        RECT 72.640 183.460 72.900 183.780 ;
        RECT 73.620 183.440 73.760 185.500 ;
        RECT 74.540 185.480 74.680 190.600 ;
        RECT 76.380 190.240 76.520 193.660 ;
        RECT 80.060 191.260 80.200 196.720 ;
        RECT 85.520 195.360 85.780 195.680 ;
        RECT 85.580 194.660 85.720 195.360 ;
        RECT 85.520 194.340 85.780 194.660 ;
        RECT 85.060 193.320 85.320 193.640 ;
        RECT 80.000 190.940 80.260 191.260 ;
        RECT 76.320 189.920 76.580 190.240 ;
        RECT 76.380 186.160 76.520 189.920 ;
        RECT 76.800 189.385 78.680 189.755 ;
        RECT 76.320 185.840 76.580 186.160 ;
        RECT 74.480 185.160 74.740 185.480 ;
        RECT 75.860 184.820 76.120 185.140 ;
        RECT 74.480 184.480 74.740 184.800 ;
        RECT 74.020 183.460 74.280 183.780 ;
        RECT 73.560 183.350 73.820 183.440 ;
        RECT 73.160 183.210 73.820 183.350 ;
        RECT 72.640 183.010 72.900 183.100 ;
        RECT 72.240 182.870 72.900 183.010 ;
        RECT 72.640 182.780 72.900 182.870 ;
        RECT 72.640 182.100 72.900 182.420 ;
        RECT 72.700 180.380 72.840 182.100 ;
        RECT 73.160 180.380 73.300 183.210 ;
        RECT 73.560 183.120 73.820 183.210 ;
        RECT 73.560 182.440 73.820 182.760 ;
        RECT 72.640 180.060 72.900 180.380 ;
        RECT 73.100 180.060 73.360 180.380 ;
        RECT 71.260 179.720 71.520 180.040 ;
        RECT 70.330 177.485 70.610 177.855 ;
        RECT 69.880 174.620 70.140 174.940 ;
        RECT 68.960 174.280 69.220 174.600 ;
        RECT 69.020 172.220 69.160 174.280 ;
        RECT 68.960 171.900 69.220 172.220 ;
        RECT 67.580 169.860 67.840 170.180 ;
        RECT 66.660 166.120 66.920 166.440 ;
        RECT 66.720 161.340 66.860 166.120 ;
        RECT 67.120 162.720 67.380 163.040 ;
        RECT 66.660 161.020 66.920 161.340 ;
        RECT 67.180 161.000 67.320 162.720 ;
        RECT 67.120 160.680 67.380 161.000 ;
        RECT 67.120 160.000 67.380 160.320 ;
        RECT 67.180 156.580 67.320 160.000 ;
        RECT 67.120 156.260 67.380 156.580 ;
        RECT 65.740 155.415 66.000 155.560 ;
        RECT 65.730 155.045 66.010 155.415 ;
        RECT 64.360 152.860 64.620 153.180 ;
        RECT 65.740 152.520 66.000 152.840 ;
        RECT 65.800 151.140 65.940 152.520 ;
        RECT 61.140 150.820 61.400 151.140 ;
        RECT 65.740 150.820 66.000 151.140 ;
        RECT 53.320 150.140 53.580 150.460 ;
        RECT 53.780 150.140 54.040 150.460 ;
        RECT 56.540 150.140 56.800 150.460 ;
        RECT 58.840 150.140 59.100 150.460 ;
        RECT 63.900 150.140 64.160 150.460 ;
        RECT 53.380 147.740 53.520 150.140 ;
        RECT 52.400 147.420 52.660 147.740 ;
        RECT 53.320 147.420 53.580 147.740 ;
        RECT 51.940 147.080 52.200 147.400 ;
        RECT 51.480 146.740 51.740 147.060 ;
        RECT 52.000 145.700 52.140 147.080 ;
        RECT 51.020 145.380 51.280 145.700 ;
        RECT 51.940 145.380 52.200 145.700 ;
        RECT 49.640 144.700 49.900 145.020 ;
        RECT 49.240 144.280 49.840 144.420 ;
        RECT 50.560 144.360 50.820 144.680 ;
        RECT 46.420 141.980 46.680 142.300 ;
        RECT 45.960 141.640 46.220 141.960 ;
        RECT 46.800 140.425 48.680 140.795 ;
        RECT 47.800 138.240 48.060 138.560 ;
        RECT 45.500 136.540 45.760 136.860 ;
        RECT 47.860 136.520 48.000 138.240 ;
        RECT 48.260 137.220 48.520 137.540 ;
        RECT 48.320 136.520 48.460 137.220 ;
        RECT 47.800 136.430 48.060 136.520 ;
        RECT 46.480 136.290 48.060 136.430 ;
        RECT 46.480 134.140 46.620 136.290 ;
        RECT 47.800 136.200 48.060 136.290 ;
        RECT 48.260 136.200 48.520 136.520 ;
        RECT 49.180 135.860 49.440 136.180 ;
        RECT 46.800 134.985 48.680 135.355 ;
        RECT 46.420 133.820 46.680 134.140 ;
        RECT 49.240 133.800 49.380 135.860 ;
        RECT 49.180 133.480 49.440 133.800 ;
        RECT 49.170 131.925 49.450 132.295 ;
        RECT 49.240 130.740 49.380 131.925 ;
        RECT 49.180 130.420 49.440 130.740 ;
        RECT 46.800 129.545 48.680 129.915 ;
        RECT 45.040 129.060 45.300 129.380 ;
        RECT 45.960 128.380 46.220 128.700 ;
        RECT 46.020 125.640 46.160 128.380 ;
        RECT 44.580 125.320 44.840 125.640 ;
        RECT 45.960 125.320 46.220 125.640 ;
        RECT 46.420 125.320 46.680 125.640 ;
        RECT 45.960 124.640 46.220 124.960 ;
        RECT 46.020 122.580 46.160 124.640 ;
        RECT 45.960 122.260 46.220 122.580 ;
        RECT 46.480 120.540 46.620 125.320 ;
        RECT 46.800 124.105 48.680 124.475 ;
        RECT 46.880 122.260 47.140 122.580 ;
        RECT 46.940 120.540 47.080 122.260 ;
        RECT 46.420 120.450 46.680 120.540 ;
        RECT 46.020 120.310 46.680 120.450 ;
        RECT 45.500 119.880 45.760 120.200 ;
        RECT 45.040 119.200 45.300 119.520 ;
        RECT 45.100 117.820 45.240 119.200 ;
        RECT 45.040 117.500 45.300 117.820 ;
        RECT 45.560 115.780 45.700 119.880 ;
        RECT 46.020 116.800 46.160 120.310 ;
        RECT 46.420 120.220 46.680 120.310 ;
        RECT 46.880 120.220 47.140 120.540 ;
        RECT 46.420 119.540 46.680 119.860 ;
        RECT 46.480 117.820 46.620 119.540 ;
        RECT 46.800 118.665 48.680 119.035 ;
        RECT 46.420 117.500 46.680 117.820 ;
        RECT 45.960 116.480 46.220 116.800 ;
        RECT 45.500 115.460 45.760 115.780 ;
        RECT 46.020 115.100 46.160 116.480 ;
        RECT 45.960 114.780 46.220 115.100 ;
        RECT 46.800 113.225 48.680 113.595 ;
        RECT 49.240 112.720 49.380 130.420 ;
        RECT 49.700 129.380 49.840 144.280 ;
        RECT 50.100 138.240 50.360 138.560 ;
        RECT 50.160 134.140 50.300 138.240 ;
        RECT 50.620 136.860 50.760 144.360 ;
        RECT 53.380 142.300 53.520 147.420 ;
        RECT 53.840 145.700 53.980 150.140 ;
        RECT 54.240 149.860 54.500 150.120 ;
        RECT 54.240 149.800 54.900 149.860 ;
        RECT 54.300 149.720 54.900 149.800 ;
        RECT 54.760 148.420 54.900 149.720 ;
        RECT 54.700 148.100 54.960 148.420 ;
        RECT 54.760 147.400 54.900 148.100 ;
        RECT 56.600 147.400 56.740 150.140 ;
        RECT 57.000 147.760 57.260 148.080 ;
        RECT 54.700 147.310 54.960 147.400 ;
        RECT 56.540 147.310 56.800 147.400 ;
        RECT 54.300 147.170 54.960 147.310 ;
        RECT 53.780 145.380 54.040 145.700 ;
        RECT 54.300 142.380 54.440 147.170 ;
        RECT 54.700 147.080 54.960 147.170 ;
        RECT 56.140 147.170 56.800 147.310 ;
        RECT 55.160 145.040 55.420 145.360 ;
        RECT 54.700 144.360 54.960 144.680 ;
        RECT 53.320 141.980 53.580 142.300 ;
        RECT 53.840 142.240 54.440 142.380 ;
        RECT 53.380 137.540 53.520 141.980 ;
        RECT 53.840 141.960 53.980 142.240 ;
        RECT 53.780 141.640 54.040 141.960 ;
        RECT 53.840 138.560 53.980 141.640 ;
        RECT 53.780 138.240 54.040 138.560 ;
        RECT 51.020 137.220 51.280 137.540 ;
        RECT 53.320 137.220 53.580 137.540 ;
        RECT 50.560 136.540 50.820 136.860 ;
        RECT 50.560 135.860 50.820 136.180 ;
        RECT 50.620 134.820 50.760 135.860 ;
        RECT 50.560 134.500 50.820 134.820 ;
        RECT 51.080 134.220 51.220 137.220 ;
        RECT 54.760 136.860 54.900 144.360 ;
        RECT 55.220 139.240 55.360 145.040 ;
        RECT 56.140 141.960 56.280 147.170 ;
        RECT 56.540 147.080 56.800 147.170 ;
        RECT 56.080 141.640 56.340 141.960 ;
        RECT 56.140 140.340 56.280 141.640 ;
        RECT 55.680 140.200 56.280 140.340 ;
        RECT 55.160 138.920 55.420 139.240 ;
        RECT 54.700 136.540 54.960 136.860 ;
        RECT 52.400 135.860 52.660 136.180 ;
        RECT 51.940 135.520 52.200 135.840 ;
        RECT 50.620 134.140 51.220 134.220 ;
        RECT 50.100 133.820 50.360 134.140 ;
        RECT 50.560 134.080 51.220 134.140 ;
        RECT 50.560 133.820 50.820 134.080 ;
        RECT 50.620 133.120 50.760 133.820 ;
        RECT 50.560 132.800 50.820 133.120 ;
        RECT 49.640 129.060 49.900 129.380 ;
        RECT 50.100 119.880 50.360 120.200 ;
        RECT 49.640 119.200 49.900 119.520 ;
        RECT 49.700 114.760 49.840 119.200 ;
        RECT 50.160 115.100 50.300 119.880 ;
        RECT 51.020 119.200 51.280 119.520 ;
        RECT 51.080 118.160 51.220 119.200 ;
        RECT 51.020 117.840 51.280 118.160 ;
        RECT 50.100 114.780 50.360 115.100 ;
        RECT 49.640 114.440 49.900 114.760 ;
        RECT 49.180 112.400 49.440 112.720 ;
        RECT 44.180 111.740 46.160 111.880 ;
        RECT 46.020 106.940 46.160 111.740 ;
        RECT 50.560 111.720 50.820 112.040 ;
        RECT 46.800 107.785 48.680 108.155 ;
        RECT 36.760 106.620 37.020 106.940 ;
        RECT 38.600 106.620 38.860 106.940 ;
        RECT 41.360 106.620 41.620 106.940 ;
        RECT 45.960 106.620 46.220 106.940 ;
        RECT 50.100 106.620 50.360 106.940 ;
        RECT 35.380 106.280 35.640 106.600 ;
        RECT 35.440 104.220 35.580 106.280 ;
        RECT 36.300 105.600 36.560 105.920 ;
        RECT 36.360 104.220 36.500 105.600 ;
        RECT 36.820 104.900 36.960 106.620 ;
        RECT 49.640 106.280 49.900 106.600 ;
        RECT 43.200 105.600 43.460 105.920 ;
        RECT 48.260 105.600 48.520 105.920 ;
        RECT 36.760 104.580 37.020 104.900 ;
        RECT 35.380 103.900 35.640 104.220 ;
        RECT 36.300 103.900 36.560 104.220 ;
        RECT 34.000 101.520 34.260 101.840 ;
        RECT 36.820 101.500 36.960 104.580 ;
        RECT 43.260 103.540 43.400 105.600 ;
        RECT 48.320 104.220 48.460 105.600 ;
        RECT 49.700 104.300 49.840 106.280 ;
        RECT 50.160 104.900 50.300 106.620 ;
        RECT 50.100 104.580 50.360 104.900 ;
        RECT 50.620 104.560 50.760 111.720 ;
        RECT 52.000 109.320 52.140 135.520 ;
        RECT 52.460 134.140 52.600 135.860 ;
        RECT 52.400 133.820 52.660 134.140 ;
        RECT 54.760 128.360 54.900 136.540 ;
        RECT 55.680 136.180 55.820 140.200 ;
        RECT 56.080 139.260 56.340 139.580 ;
        RECT 55.620 135.860 55.880 136.180 ;
        RECT 56.140 134.480 56.280 139.260 ;
        RECT 56.540 135.520 56.800 135.840 ;
        RECT 56.600 134.820 56.740 135.520 ;
        RECT 56.540 134.500 56.800 134.820 ;
        RECT 56.080 134.160 56.340 134.480 ;
        RECT 55.620 133.140 55.880 133.460 ;
        RECT 55.680 129.380 55.820 133.140 ;
        RECT 56.600 129.380 56.740 134.500 ;
        RECT 55.620 129.060 55.880 129.380 ;
        RECT 56.540 129.060 56.800 129.380 ;
        RECT 54.700 128.040 54.960 128.360 ;
        RECT 54.760 125.980 54.900 128.040 ;
        RECT 55.680 126.320 55.820 129.060 ;
        RECT 55.620 126.000 55.880 126.320 ;
        RECT 54.700 125.660 54.960 125.980 ;
        RECT 55.680 123.940 55.820 126.000 ;
        RECT 55.620 123.620 55.880 123.940 ;
        RECT 54.700 117.500 54.960 117.820 ;
        RECT 54.760 115.780 54.900 117.500 ;
        RECT 56.540 117.160 56.800 117.480 ;
        RECT 54.700 115.460 54.960 115.780 ;
        RECT 51.940 109.000 52.200 109.320 ;
        RECT 55.620 108.320 55.880 108.640 ;
        RECT 55.680 107.280 55.820 108.320 ;
        RECT 55.620 106.960 55.880 107.280 ;
        RECT 52.400 106.280 52.660 106.600 ;
        RECT 56.600 106.510 56.740 117.160 ;
        RECT 57.060 109.320 57.200 147.760 ;
        RECT 58.900 147.060 59.040 150.140 ;
        RECT 60.220 149.460 60.480 149.780 ;
        RECT 58.840 146.740 59.100 147.060 ;
        RECT 59.300 146.400 59.560 146.720 ;
        RECT 59.360 145.360 59.500 146.400 ;
        RECT 59.300 145.040 59.560 145.360 ;
        RECT 58.840 143.680 59.100 144.000 ;
        RECT 58.900 141.620 59.040 143.680 ;
        RECT 59.360 142.980 59.500 145.040 ;
        RECT 59.300 142.660 59.560 142.980 ;
        RECT 58.840 141.300 59.100 141.620 ;
        RECT 59.760 135.520 60.020 135.840 ;
        RECT 59.820 134.140 59.960 135.520 ;
        RECT 59.760 133.820 60.020 134.140 ;
        RECT 60.280 133.540 60.420 149.460 ;
        RECT 61.800 148.585 63.680 148.955 ;
        RECT 63.960 146.720 64.100 150.140 ;
        RECT 65.740 149.800 66.000 150.120 ;
        RECT 64.820 149.460 65.080 149.780 ;
        RECT 64.880 147.740 65.020 149.460 ;
        RECT 65.280 149.120 65.540 149.440 ;
        RECT 64.820 147.420 65.080 147.740 ;
        RECT 63.900 146.400 64.160 146.720 ;
        RECT 64.880 144.680 65.020 147.420 ;
        RECT 64.820 144.360 65.080 144.680 ;
        RECT 63.900 144.020 64.160 144.340 ;
        RECT 61.800 143.145 63.680 143.515 ;
        RECT 63.960 141.280 64.100 144.020 ;
        RECT 63.900 140.960 64.160 141.280 ;
        RECT 61.140 139.940 61.400 140.260 ;
        RECT 60.680 139.260 60.940 139.580 ;
        RECT 60.740 137.540 60.880 139.260 ;
        RECT 60.680 137.220 60.940 137.540 ;
        RECT 60.680 135.860 60.940 136.180 ;
        RECT 59.820 133.400 60.420 133.540 ;
        RECT 57.920 127.360 58.180 127.680 ;
        RECT 57.980 125.640 58.120 127.360 ;
        RECT 57.920 125.320 58.180 125.640 ;
        RECT 57.460 123.280 57.720 123.600 ;
        RECT 57.520 121.220 57.660 123.280 ;
        RECT 59.820 122.660 59.960 133.400 ;
        RECT 60.740 125.640 60.880 135.860 ;
        RECT 61.200 135.840 61.340 139.940 ;
        RECT 61.800 137.705 63.680 138.075 ;
        RECT 61.140 135.520 61.400 135.840 ;
        RECT 63.960 134.140 64.100 140.960 ;
        RECT 65.340 139.580 65.480 149.120 ;
        RECT 65.800 147.400 65.940 149.800 ;
        RECT 65.740 147.080 66.000 147.400 ;
        RECT 65.740 144.700 66.000 145.020 ;
        RECT 65.800 140.260 65.940 144.700 ;
        RECT 65.740 139.940 66.000 140.260 ;
        RECT 65.280 139.260 65.540 139.580 ;
        RECT 64.360 138.580 64.620 138.900 ;
        RECT 64.420 136.520 64.560 138.580 ;
        RECT 65.340 137.540 65.480 139.260 ;
        RECT 65.280 137.220 65.540 137.540 ;
        RECT 65.340 136.940 65.480 137.220 ;
        RECT 64.880 136.800 65.480 136.940 ;
        RECT 65.800 136.860 65.940 139.940 ;
        RECT 66.200 139.260 66.460 139.580 ;
        RECT 64.360 136.200 64.620 136.520 ;
        RECT 64.420 134.480 64.560 136.200 ;
        RECT 64.360 134.160 64.620 134.480 ;
        RECT 64.880 134.140 65.020 136.800 ;
        RECT 65.740 136.540 66.000 136.860 ;
        RECT 65.280 135.860 65.540 136.180 ;
        RECT 65.340 134.140 65.480 135.860 ;
        RECT 63.900 133.820 64.160 134.140 ;
        RECT 64.820 133.820 65.080 134.140 ;
        RECT 65.280 133.820 65.540 134.140 ;
        RECT 65.740 133.820 66.000 134.140 ;
        RECT 61.800 132.265 63.680 132.635 ;
        RECT 63.960 129.040 64.100 133.820 ;
        RECT 64.820 131.100 65.080 131.420 ;
        RECT 64.360 130.420 64.620 130.740 ;
        RECT 63.900 128.720 64.160 129.040 ;
        RECT 63.960 128.360 64.100 128.720 ;
        RECT 63.900 128.040 64.160 128.360 ;
        RECT 61.800 126.825 63.680 127.195 ;
        RECT 60.680 125.320 60.940 125.640 ;
        RECT 60.220 124.640 60.480 124.960 ;
        RECT 60.280 123.260 60.420 124.640 ;
        RECT 60.740 123.940 60.880 125.320 ;
        RECT 60.680 123.620 60.940 123.940 ;
        RECT 60.220 122.940 60.480 123.260 ;
        RECT 59.820 122.520 60.420 122.660 ;
        RECT 57.460 120.900 57.720 121.220 ;
        RECT 57.920 119.880 58.180 120.200 ;
        RECT 57.980 117.820 58.120 119.880 ;
        RECT 57.920 117.500 58.180 117.820 ;
        RECT 59.760 117.500 60.020 117.820 ;
        RECT 59.820 109.320 59.960 117.500 ;
        RECT 60.280 111.880 60.420 122.520 ;
        RECT 60.740 121.220 60.880 123.620 ;
        RECT 63.960 123.260 64.100 128.040 ;
        RECT 64.420 123.260 64.560 130.420 ;
        RECT 63.900 122.940 64.160 123.260 ;
        RECT 64.360 122.940 64.620 123.260 ;
        RECT 61.800 121.385 63.680 121.755 ;
        RECT 60.680 120.900 60.940 121.220 ;
        RECT 62.060 119.540 62.320 119.860 ;
        RECT 62.120 118.500 62.260 119.540 ;
        RECT 64.420 118.500 64.560 122.940 ;
        RECT 64.880 122.920 65.020 131.100 ;
        RECT 65.800 130.740 65.940 133.820 ;
        RECT 65.740 130.420 66.000 130.740 ;
        RECT 66.260 130.400 66.400 139.260 ;
        RECT 67.640 138.900 67.780 169.860 ;
        RECT 68.500 166.460 68.760 166.780 ;
        RECT 68.560 163.720 68.700 166.460 ;
        RECT 69.020 165.760 69.160 171.900 ;
        RECT 70.400 169.160 70.540 177.485 ;
        RECT 70.800 173.600 71.060 173.920 ;
        RECT 70.860 170.180 71.000 173.600 ;
        RECT 70.800 169.860 71.060 170.180 ;
        RECT 70.340 168.840 70.600 169.160 ;
        RECT 70.400 167.460 70.540 168.840 ;
        RECT 70.340 167.140 70.600 167.460 ;
        RECT 68.960 165.440 69.220 165.760 ;
        RECT 68.500 163.400 68.760 163.720 ;
        RECT 68.030 158.445 68.310 158.815 ;
        RECT 68.100 152.695 68.240 158.445 ;
        RECT 68.030 152.325 68.310 152.695 ;
        RECT 68.500 152.520 68.760 152.840 ;
        RECT 68.100 139.580 68.240 152.325 ;
        RECT 68.560 142.300 68.700 152.520 ;
        RECT 69.020 144.340 69.160 165.440 ;
        RECT 69.880 160.000 70.140 160.320 ;
        RECT 69.420 157.960 69.680 158.280 ;
        RECT 69.480 153.180 69.620 157.960 ;
        RECT 69.940 154.880 70.080 160.000 ;
        RECT 70.400 158.280 70.540 167.140 ;
        RECT 71.320 166.860 71.460 179.720 ;
        RECT 73.100 179.380 73.360 179.700 ;
        RECT 73.160 178.340 73.300 179.380 ;
        RECT 71.720 178.020 71.980 178.340 ;
        RECT 73.100 178.020 73.360 178.340 ;
        RECT 71.780 177.175 71.920 178.020 ;
        RECT 72.630 177.485 72.910 177.855 ;
        RECT 72.640 177.340 72.900 177.485 ;
        RECT 71.710 176.805 71.990 177.175 ;
        RECT 72.700 174.600 72.840 177.340 ;
        RECT 72.640 174.280 72.900 174.600 ;
        RECT 73.620 171.620 73.760 182.440 ;
        RECT 74.080 180.040 74.220 183.460 ;
        RECT 74.020 179.720 74.280 180.040 ;
        RECT 74.020 177.340 74.280 177.660 ;
        RECT 70.860 166.780 71.460 166.860 ;
        RECT 70.800 166.720 71.460 166.780 ;
        RECT 70.800 166.460 71.060 166.720 ;
        RECT 71.320 161.340 71.460 166.720 ;
        RECT 72.700 171.480 73.760 171.620 ;
        RECT 71.260 161.020 71.520 161.340 ;
        RECT 70.800 160.340 71.060 160.660 ;
        RECT 70.860 158.960 71.000 160.340 ;
        RECT 71.720 158.980 71.980 159.300 ;
        RECT 70.800 158.640 71.060 158.960 ;
        RECT 71.780 158.815 71.920 158.980 ;
        RECT 71.710 158.445 71.990 158.815 ;
        RECT 70.340 157.960 70.600 158.280 ;
        RECT 69.880 154.560 70.140 154.880 ;
        RECT 69.940 153.520 70.080 154.560 ;
        RECT 70.340 153.540 70.600 153.860 ;
        RECT 69.880 153.200 70.140 153.520 ;
        RECT 69.420 152.860 69.680 153.180 ;
        RECT 69.480 150.460 69.620 152.860 ;
        RECT 70.400 152.160 70.540 153.540 ;
        RECT 70.800 152.580 71.060 152.840 ;
        RECT 71.720 152.580 71.980 152.840 ;
        RECT 70.800 152.520 71.980 152.580 ;
        RECT 70.860 152.440 71.920 152.520 ;
        RECT 70.340 151.840 70.600 152.160 ;
        RECT 69.420 150.140 69.680 150.460 ;
        RECT 69.420 144.360 69.680 144.680 ;
        RECT 68.960 144.020 69.220 144.340 ;
        RECT 68.960 142.320 69.220 142.640 ;
        RECT 68.500 141.980 68.760 142.300 ;
        RECT 68.560 141.280 68.700 141.980 ;
        RECT 68.500 140.960 68.760 141.280 ;
        RECT 68.040 139.260 68.300 139.580 ;
        RECT 67.580 138.580 67.840 138.900 ;
        RECT 66.660 138.240 66.920 138.560 ;
        RECT 66.720 136.180 66.860 138.240 ;
        RECT 66.660 135.860 66.920 136.180 ;
        RECT 68.040 130.420 68.300 130.740 ;
        RECT 66.200 130.080 66.460 130.400 ;
        RECT 66.260 129.380 66.400 130.080 ;
        RECT 66.200 129.060 66.460 129.380 ;
        RECT 68.100 128.700 68.240 130.420 ;
        RECT 68.500 128.720 68.760 129.040 ;
        RECT 68.040 128.380 68.300 128.700 ;
        RECT 68.560 125.640 68.700 128.720 ;
        RECT 68.500 125.320 68.760 125.640 ;
        RECT 64.820 122.600 65.080 122.920 ;
        RECT 68.040 121.920 68.300 122.240 ;
        RECT 62.060 118.180 62.320 118.500 ;
        RECT 64.360 118.180 64.620 118.500 ;
        RECT 66.660 117.840 66.920 118.160 ;
        RECT 61.800 115.945 63.680 116.315 ;
        RECT 66.720 115.780 66.860 117.840 ;
        RECT 66.660 115.460 66.920 115.780 ;
        RECT 68.100 114.760 68.240 121.920 ;
        RECT 68.040 114.440 68.300 114.760 ;
        RECT 60.280 111.740 60.880 111.880 ;
        RECT 57.000 109.000 57.260 109.320 ;
        RECT 59.760 109.000 60.020 109.320 ;
        RECT 60.220 109.000 60.480 109.320 ;
        RECT 57.920 108.320 58.180 108.640 ;
        RECT 57.000 106.510 57.260 106.600 ;
        RECT 56.600 106.370 57.260 106.510 ;
        RECT 48.260 103.900 48.520 104.220 ;
        RECT 49.700 104.160 50.300 104.300 ;
        RECT 50.560 104.240 50.820 104.560 ;
        RECT 39.060 103.220 39.320 103.540 ;
        RECT 43.200 103.220 43.460 103.540 ;
        RECT 36.760 101.180 37.020 101.500 ;
        RECT 31.800 99.625 33.680 99.995 ;
        RECT 31.780 88.660 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 30.380 88.520 33.000 88.660 ;
        RECT 31.780 85.510 33.000 88.520 ;
        RECT 37.680 88.660 38.970 88.780 ;
        RECT 39.120 88.660 39.260 103.220 ;
        RECT 44.120 102.880 44.380 103.200 ;
        RECT 44.180 89.530 44.320 102.880 ;
        RECT 46.800 102.345 48.680 102.715 ;
        RECT 37.680 88.520 39.260 88.660 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 50.160 89.210 50.300 104.160 ;
        RECT 52.460 103.880 52.600 106.280 ;
        RECT 56.600 104.900 56.740 106.370 ;
        RECT 57.000 106.280 57.260 106.370 ;
        RECT 57.000 105.600 57.260 105.920 ;
        RECT 56.540 104.580 56.800 104.900 ;
        RECT 57.060 104.300 57.200 105.600 ;
        RECT 56.600 104.160 57.200 104.300 ;
        RECT 57.980 104.220 58.120 108.320 ;
        RECT 60.280 106.940 60.420 109.000 ;
        RECT 60.740 106.940 60.880 111.740 ;
        RECT 61.800 110.505 63.680 110.875 ;
        RECT 69.020 109.320 69.160 142.320 ;
        RECT 69.480 136.520 69.620 144.360 ;
        RECT 69.880 143.680 70.140 144.000 ;
        RECT 69.940 141.960 70.080 143.680 ;
        RECT 69.880 141.640 70.140 141.960 ;
        RECT 70.400 139.240 70.540 151.840 ;
        RECT 70.860 150.460 71.000 152.440 ;
        RECT 72.180 152.180 72.440 152.500 ;
        RECT 70.800 150.140 71.060 150.460 ;
        RECT 70.860 147.740 71.000 150.140 ;
        RECT 70.800 147.420 71.060 147.740 ;
        RECT 72.240 147.400 72.380 152.180 ;
        RECT 72.180 147.080 72.440 147.400 ;
        RECT 70.800 144.020 71.060 144.340 ;
        RECT 70.860 141.960 71.000 144.020 ;
        RECT 70.800 141.640 71.060 141.960 ;
        RECT 70.340 138.920 70.600 139.240 ;
        RECT 69.420 136.200 69.680 136.520 ;
        RECT 69.480 131.420 69.620 136.200 ;
        RECT 69.420 131.100 69.680 131.420 ;
        RECT 70.860 130.820 71.000 141.640 ;
        RECT 72.180 140.960 72.440 141.280 ;
        RECT 72.240 139.920 72.380 140.960 ;
        RECT 72.180 139.600 72.440 139.920 ;
        RECT 72.700 131.080 72.840 171.480 ;
        RECT 74.080 166.440 74.220 177.340 ;
        RECT 74.020 166.120 74.280 166.440 ;
        RECT 73.100 165.440 73.360 165.760 ;
        RECT 73.160 163.720 73.300 165.440 ;
        RECT 73.100 163.400 73.360 163.720 ;
        RECT 73.160 158.280 73.300 163.400 ;
        RECT 74.540 161.250 74.680 184.480 ;
        RECT 75.920 183.100 76.060 184.820 ;
        RECT 75.860 182.780 76.120 183.100 ;
        RECT 75.920 182.420 76.060 182.780 ;
        RECT 75.860 182.100 76.120 182.420 ;
        RECT 74.940 181.760 75.200 182.080 ;
        RECT 76.380 181.820 76.520 185.840 ;
        RECT 85.120 185.820 85.260 193.320 ;
        RECT 85.580 191.940 85.720 194.340 ;
        RECT 86.960 194.320 87.100 199.100 ;
        RECT 91.800 197.545 93.680 197.915 ;
        RECT 93.800 196.380 94.060 196.700 ;
        RECT 90.120 195.700 90.380 196.020 ;
        RECT 90.180 194.660 90.320 195.700 ;
        RECT 90.120 194.340 90.380 194.660 ;
        RECT 86.900 194.000 87.160 194.320 ;
        RECT 85.980 193.660 86.240 193.980 ;
        RECT 90.120 193.660 90.380 193.980 ;
        RECT 85.520 191.620 85.780 191.940 ;
        RECT 85.060 185.500 85.320 185.820 ;
        RECT 76.800 183.945 78.680 184.315 ;
        RECT 76.780 182.780 77.040 183.100 ;
        RECT 76.840 181.820 76.980 182.780 ;
        RECT 85.120 182.080 85.260 185.500 ;
        RECT 75.000 177.660 75.140 181.760 ;
        RECT 75.920 181.680 76.980 181.820 ;
        RECT 79.540 181.760 79.800 182.080 ;
        RECT 85.060 181.760 85.320 182.080 ;
        RECT 75.920 180.380 76.060 181.680 ;
        RECT 79.080 180.400 79.340 180.720 ;
        RECT 75.860 180.060 76.120 180.380 ;
        RECT 76.320 179.720 76.580 180.040 ;
        RECT 76.380 177.660 76.520 179.720 ;
        RECT 78.610 179.525 78.890 179.895 ;
        RECT 78.680 179.360 78.820 179.525 ;
        RECT 78.620 179.040 78.880 179.360 ;
        RECT 76.800 178.505 78.680 178.875 ;
        RECT 74.940 177.340 75.200 177.660 ;
        RECT 76.320 177.340 76.580 177.660 ;
        RECT 77.700 177.340 77.960 177.660 ;
        RECT 78.160 177.340 78.420 177.660 ;
        RECT 75.000 176.640 75.140 177.340 ;
        RECT 74.940 176.320 75.200 176.640 ;
        RECT 76.380 175.280 76.520 177.340 ;
        RECT 77.760 175.620 77.900 177.340 ;
        RECT 78.220 177.175 78.360 177.340 ;
        RECT 79.140 177.320 79.280 180.400 ;
        RECT 79.600 180.380 79.740 181.760 ;
        RECT 82.300 180.740 82.560 181.060 ;
        RECT 79.540 180.060 79.800 180.380 ;
        RECT 81.380 179.720 81.640 180.040 ;
        RECT 81.840 179.720 82.100 180.040 ;
        RECT 79.540 177.680 79.800 178.000 ;
        RECT 78.150 176.805 78.430 177.175 ;
        RECT 79.080 177.000 79.340 177.320 ;
        RECT 77.700 175.300 77.960 175.620 ;
        RECT 76.320 174.960 76.580 175.280 ;
        RECT 78.220 174.600 78.360 176.805 ;
        RECT 78.160 174.280 78.420 174.600 ;
        RECT 76.800 173.065 78.680 173.435 ;
        RECT 76.320 168.160 76.580 168.480 ;
        RECT 79.080 168.160 79.340 168.480 ;
        RECT 74.940 166.120 75.200 166.440 ;
        RECT 73.620 161.110 74.680 161.250 ;
        RECT 73.100 157.960 73.360 158.280 ;
        RECT 73.090 156.405 73.370 156.775 ;
        RECT 69.940 130.680 71.000 130.820 ;
        RECT 72.640 130.760 72.900 131.080 ;
        RECT 69.940 125.640 70.080 130.680 ;
        RECT 70.340 130.080 70.600 130.400 ;
        RECT 71.720 130.080 71.980 130.400 ;
        RECT 70.400 125.640 70.540 130.080 ;
        RECT 71.780 125.640 71.920 130.080 ;
        RECT 72.180 128.380 72.440 128.700 ;
        RECT 72.240 126.660 72.380 128.380 ;
        RECT 72.180 126.340 72.440 126.660 ;
        RECT 69.880 125.550 70.140 125.640 ;
        RECT 69.480 125.410 70.140 125.550 ;
        RECT 69.480 117.480 69.620 125.410 ;
        RECT 69.880 125.320 70.140 125.410 ;
        RECT 70.340 125.320 70.600 125.640 ;
        RECT 71.720 125.320 71.980 125.640 ;
        RECT 69.880 124.640 70.140 124.960 ;
        RECT 69.940 120.200 70.080 124.640 ;
        RECT 73.160 123.260 73.300 156.405 ;
        RECT 73.620 153.860 73.760 161.110 ;
        RECT 74.020 160.000 74.280 160.320 ;
        RECT 74.080 158.280 74.220 160.000 ;
        RECT 74.020 157.960 74.280 158.280 ;
        RECT 74.080 157.600 74.220 157.960 ;
        RECT 74.020 157.280 74.280 157.600 ;
        RECT 74.080 156.240 74.220 157.280 ;
        RECT 74.020 155.920 74.280 156.240 ;
        RECT 74.480 155.580 74.740 155.900 ;
        RECT 74.540 155.415 74.680 155.580 ;
        RECT 74.470 155.045 74.750 155.415 ;
        RECT 73.560 153.540 73.820 153.860 ;
        RECT 73.620 152.500 73.760 153.540 ;
        RECT 74.020 153.090 74.280 153.180 ;
        RECT 75.000 153.090 75.140 166.120 ;
        RECT 75.400 163.060 75.660 163.380 ;
        RECT 75.460 156.775 75.600 163.060 ;
        RECT 76.380 158.620 76.520 168.160 ;
        RECT 76.800 167.625 78.680 167.995 ;
        RECT 78.620 165.780 78.880 166.100 ;
        RECT 78.680 164.060 78.820 165.780 ;
        RECT 78.620 163.740 78.880 164.060 ;
        RECT 79.140 163.380 79.280 168.160 ;
        RECT 79.080 163.060 79.340 163.380 ;
        RECT 76.800 162.185 78.680 162.555 ;
        RECT 76.320 158.300 76.580 158.620 ;
        RECT 79.080 157.960 79.340 158.280 ;
        RECT 76.320 157.620 76.580 157.940 ;
        RECT 75.860 157.280 76.120 157.600 ;
        RECT 75.390 156.405 75.670 156.775 ;
        RECT 74.020 152.950 75.140 153.090 ;
        RECT 74.020 152.860 74.280 152.950 ;
        RECT 73.560 152.180 73.820 152.500 ;
        RECT 73.560 148.100 73.820 148.420 ;
        RECT 73.620 146.720 73.760 148.100 ;
        RECT 73.560 146.400 73.820 146.720 ;
        RECT 74.080 136.860 74.220 152.860 ;
        RECT 74.940 151.840 75.200 152.160 ;
        RECT 75.000 150.800 75.140 151.840 ;
        RECT 74.940 150.480 75.200 150.800 ;
        RECT 75.920 150.460 76.060 157.280 ;
        RECT 76.380 155.560 76.520 157.620 ;
        RECT 76.800 156.745 78.680 157.115 ;
        RECT 79.140 156.490 79.280 157.960 ;
        RECT 78.220 156.350 79.280 156.490 ;
        RECT 78.220 155.900 78.360 156.350 ;
        RECT 78.160 155.580 78.420 155.900 ;
        RECT 78.620 155.580 78.880 155.900 ;
        RECT 76.320 155.240 76.580 155.560 ;
        RECT 78.680 155.220 78.820 155.580 ;
        RECT 78.620 154.900 78.880 155.220 ;
        RECT 76.320 154.560 76.580 154.880 ;
        RECT 75.860 150.140 76.120 150.460 ;
        RECT 75.860 149.120 76.120 149.440 ;
        RECT 75.400 144.020 75.660 144.340 ;
        RECT 74.940 138.920 75.200 139.240 ;
        RECT 75.000 137.540 75.140 138.920 ;
        RECT 74.940 137.220 75.200 137.540 ;
        RECT 74.480 136.880 74.740 137.200 ;
        RECT 74.020 136.540 74.280 136.860 ;
        RECT 74.080 131.420 74.220 136.540 ;
        RECT 74.540 134.820 74.680 136.880 ;
        RECT 74.480 134.500 74.740 134.820 ;
        RECT 74.020 131.100 74.280 131.420 ;
        RECT 73.100 122.940 73.360 123.260 ;
        RECT 73.160 120.200 73.300 122.940 ;
        RECT 69.880 119.880 70.140 120.200 ;
        RECT 73.100 119.880 73.360 120.200 ;
        RECT 70.800 119.540 71.060 119.860 ;
        RECT 70.860 118.580 71.000 119.540 ;
        RECT 70.860 118.440 71.460 118.580 ;
        RECT 71.320 117.480 71.460 118.440 ;
        RECT 69.420 117.160 69.680 117.480 ;
        RECT 70.800 117.160 71.060 117.480 ;
        RECT 71.260 117.160 71.520 117.480 ;
        RECT 69.480 115.100 69.620 117.160 ;
        RECT 70.860 115.780 71.000 117.160 ;
        RECT 71.320 115.780 71.460 117.160 ;
        RECT 70.800 115.460 71.060 115.780 ;
        RECT 71.260 115.460 71.520 115.780 ;
        RECT 73.560 115.460 73.820 115.780 ;
        RECT 69.420 114.780 69.680 115.100 ;
        RECT 68.960 109.000 69.220 109.320 ;
        RECT 65.280 108.320 65.540 108.640 ;
        RECT 72.180 108.320 72.440 108.640 ;
        RECT 65.340 107.280 65.480 108.320 ;
        RECT 72.240 107.280 72.380 108.320 ;
        RECT 65.280 106.960 65.540 107.280 ;
        RECT 72.180 106.960 72.440 107.280 ;
        RECT 60.220 106.620 60.480 106.940 ;
        RECT 60.680 106.620 60.940 106.940 ;
        RECT 73.620 106.600 73.760 115.460 ;
        RECT 74.080 110.340 74.220 131.100 ;
        RECT 74.940 130.080 75.200 130.400 ;
        RECT 75.000 128.700 75.140 130.080 ;
        RECT 74.940 128.380 75.200 128.700 ;
        RECT 75.460 128.100 75.600 144.020 ;
        RECT 75.000 127.960 75.600 128.100 ;
        RECT 74.020 110.020 74.280 110.340 ;
        RECT 75.000 106.940 75.140 127.960 ;
        RECT 75.400 119.200 75.660 119.520 ;
        RECT 75.460 118.160 75.600 119.200 ;
        RECT 75.400 117.840 75.660 118.160 ;
        RECT 75.920 108.980 76.060 149.120 ;
        RECT 76.380 136.520 76.520 154.560 ;
        RECT 76.800 151.305 78.680 151.675 ;
        RECT 79.600 150.120 79.740 177.680 ;
        RECT 81.440 177.570 81.580 179.720 ;
        RECT 81.900 178.340 82.040 179.720 ;
        RECT 82.360 178.340 82.500 180.740 ;
        RECT 85.120 180.380 85.260 181.760 ;
        RECT 85.580 180.720 85.720 191.620 ;
        RECT 86.040 190.240 86.180 193.660 ;
        RECT 87.820 190.260 88.080 190.580 ;
        RECT 85.980 189.920 86.240 190.240 ;
        RECT 86.040 184.800 86.180 189.920 ;
        RECT 87.880 189.220 88.020 190.260 ;
        RECT 87.820 188.900 88.080 189.220 ;
        RECT 89.200 188.220 89.460 188.540 ;
        RECT 89.260 186.500 89.400 188.220 ;
        RECT 90.180 188.200 90.320 193.660 ;
        RECT 91.040 192.640 91.300 192.960 ;
        RECT 91.100 190.920 91.240 192.640 ;
        RECT 91.800 192.105 93.680 192.475 ;
        RECT 93.860 191.940 94.000 196.380 ;
        RECT 96.620 196.360 96.760 201.480 ;
        RECT 106.800 200.265 108.680 200.635 ;
        RECT 97.940 199.440 98.200 199.760 ;
        RECT 96.560 196.040 96.820 196.360 ;
        RECT 96.620 194.320 96.760 196.040 ;
        RECT 98.000 194.660 98.140 199.440 ;
        RECT 104.380 198.760 104.640 199.080 ;
        RECT 105.760 198.760 106.020 199.080 ;
        RECT 98.400 198.080 98.660 198.400 ;
        RECT 98.460 196.360 98.600 198.080 ;
        RECT 98.400 196.040 98.660 196.360 ;
        RECT 97.940 194.340 98.200 194.660 ;
        RECT 96.560 194.000 96.820 194.320 ;
        RECT 94.720 193.660 94.980 193.980 ;
        RECT 93.800 191.620 94.060 191.940 ;
        RECT 93.800 190.940 94.060 191.260 ;
        RECT 90.580 190.600 90.840 190.920 ;
        RECT 91.040 190.600 91.300 190.920 ;
        RECT 90.640 189.220 90.780 190.600 ;
        RECT 90.580 188.900 90.840 189.220 ;
        RECT 90.120 187.880 90.380 188.200 ;
        RECT 91.040 187.880 91.300 188.200 ;
        RECT 89.200 186.180 89.460 186.500 ;
        RECT 91.100 186.160 91.240 187.880 ;
        RECT 91.800 186.665 93.680 187.035 ;
        RECT 91.040 185.840 91.300 186.160 ;
        RECT 85.980 184.480 86.240 184.800 ;
        RECT 86.440 184.480 86.700 184.800 ;
        RECT 85.520 180.400 85.780 180.720 ;
        RECT 85.060 180.060 85.320 180.380 ;
        RECT 85.120 179.895 85.260 180.060 ;
        RECT 85.050 179.525 85.330 179.895 ;
        RECT 82.760 179.040 83.020 179.360 ;
        RECT 83.680 179.040 83.940 179.360 ;
        RECT 81.840 178.020 82.100 178.340 ;
        RECT 82.300 178.020 82.560 178.340 ;
        RECT 82.820 177.660 82.960 179.040 ;
        RECT 81.840 177.570 82.100 177.660 ;
        RECT 81.440 177.430 82.100 177.570 ;
        RECT 81.840 177.340 82.100 177.430 ;
        RECT 82.760 177.340 83.020 177.660 ;
        RECT 80.460 177.000 80.720 177.320 ;
        RECT 80.000 169.180 80.260 169.500 ;
        RECT 80.060 165.760 80.200 169.180 ;
        RECT 80.000 165.440 80.260 165.760 ;
        RECT 80.060 161.000 80.200 165.440 ;
        RECT 80.000 160.680 80.260 161.000 ;
        RECT 79.990 159.125 80.270 159.495 ;
        RECT 80.000 158.980 80.260 159.125 ;
        RECT 80.520 155.300 80.660 177.000 ;
        RECT 81.900 175.620 82.040 177.340 ;
        RECT 81.840 175.300 82.100 175.620 ;
        RECT 81.840 173.940 82.100 174.260 ;
        RECT 80.920 162.720 81.180 163.040 ;
        RECT 81.900 162.780 82.040 173.940 ;
        RECT 83.220 168.160 83.480 168.480 ;
        RECT 82.760 166.120 83.020 166.440 ;
        RECT 82.820 164.740 82.960 166.120 ;
        RECT 82.760 164.420 83.020 164.740 ;
        RECT 83.280 163.720 83.420 168.160 ;
        RECT 83.740 166.180 83.880 179.040 ;
        RECT 86.040 178.000 86.180 184.480 ;
        RECT 86.500 179.700 86.640 184.480 ;
        RECT 91.100 183.100 91.240 185.840 ;
        RECT 91.040 182.780 91.300 183.100 ;
        RECT 89.660 182.100 89.920 182.420 ;
        RECT 89.720 181.060 89.860 182.100 ;
        RECT 89.660 180.740 89.920 181.060 ;
        RECT 91.100 180.040 91.240 182.780 ;
        RECT 93.860 182.760 94.000 190.940 ;
        RECT 94.780 188.055 94.920 193.660 ;
        RECT 96.620 190.920 96.760 194.000 ;
        RECT 97.940 190.940 98.200 191.260 ;
        RECT 96.560 190.600 96.820 190.920 ;
        RECT 94.710 187.685 94.990 188.055 ;
        RECT 97.480 184.480 97.740 184.800 ;
        RECT 97.540 183.780 97.680 184.480 ;
        RECT 97.480 183.460 97.740 183.780 ;
        RECT 96.100 182.780 96.360 183.100 ;
        RECT 93.800 182.440 94.060 182.760 ;
        RECT 91.800 181.225 93.680 181.595 ;
        RECT 90.580 179.720 90.840 180.040 ;
        RECT 91.040 179.720 91.300 180.040 ;
        RECT 86.440 179.380 86.700 179.700 ;
        RECT 87.360 179.040 87.620 179.360 ;
        RECT 89.200 179.040 89.460 179.360 ;
        RECT 85.980 177.680 86.240 178.000 ;
        RECT 84.140 177.340 84.400 177.660 ;
        RECT 84.200 174.600 84.340 177.340 ;
        RECT 87.420 174.940 87.560 179.040 ;
        RECT 89.260 177.660 89.400 179.040 ;
        RECT 90.640 178.340 90.780 179.720 ;
        RECT 90.580 178.020 90.840 178.340 ;
        RECT 89.200 177.340 89.460 177.660 ;
        RECT 87.360 174.620 87.620 174.940 ;
        RECT 84.140 174.280 84.400 174.600 ;
        RECT 91.100 172.900 91.240 179.720 ;
        RECT 96.160 179.360 96.300 182.780 ;
        RECT 98.000 182.760 98.140 190.940 ;
        RECT 97.940 182.440 98.200 182.760 ;
        RECT 98.460 182.420 98.600 196.040 ;
        RECT 101.160 195.360 101.420 195.680 ;
        RECT 101.220 191.260 101.360 195.360 ;
        RECT 104.440 191.940 104.580 198.760 ;
        RECT 105.820 194.320 105.960 198.760 ;
        RECT 121.800 197.545 123.680 197.915 ;
        RECT 115.420 195.700 115.680 196.020 ;
        RECT 117.720 195.700 117.980 196.020 ;
        RECT 118.180 195.700 118.440 196.020 ;
        RECT 108.980 195.360 109.240 195.680 ;
        RECT 106.800 194.825 108.680 195.195 ;
        RECT 105.760 194.000 106.020 194.320 ;
        RECT 108.060 193.320 108.320 193.640 ;
        RECT 104.380 191.620 104.640 191.940 ;
        RECT 108.120 191.600 108.260 193.320 ;
        RECT 108.060 191.280 108.320 191.600 ;
        RECT 101.160 190.940 101.420 191.260 ;
        RECT 106.220 190.940 106.480 191.260 ;
        RECT 106.280 189.220 106.420 190.940 ;
        RECT 106.800 189.385 108.680 189.755 ;
        RECT 106.220 188.900 106.480 189.220 ;
        RECT 100.240 188.560 100.500 188.880 ;
        RECT 99.320 187.200 99.580 187.520 ;
        RECT 99.780 187.200 100.040 187.520 ;
        RECT 99.380 185.820 99.520 187.200 ;
        RECT 99.840 186.500 99.980 187.200 ;
        RECT 100.300 186.500 100.440 188.560 ;
        RECT 99.780 186.180 100.040 186.500 ;
        RECT 100.240 186.180 100.500 186.500 ;
        RECT 109.040 185.820 109.180 195.360 ;
        RECT 115.480 194.660 115.620 195.700 ;
        RECT 112.660 194.340 112.920 194.660 ;
        RECT 115.420 194.340 115.680 194.660 ;
        RECT 110.820 193.320 111.080 193.640 ;
        RECT 109.440 192.640 109.700 192.960 ;
        RECT 109.500 190.580 109.640 192.640 ;
        RECT 109.900 190.940 110.160 191.260 ;
        RECT 109.440 190.260 109.700 190.580 ;
        RECT 109.960 188.540 110.100 190.940 ;
        RECT 109.900 188.220 110.160 188.540 ;
        RECT 99.320 185.500 99.580 185.820 ;
        RECT 105.300 185.500 105.560 185.820 ;
        RECT 108.980 185.500 109.240 185.820 ;
        RECT 99.380 183.100 99.520 185.500 ;
        RECT 99.320 182.780 99.580 183.100 ;
        RECT 98.400 182.100 98.660 182.420 ;
        RECT 96.100 179.040 96.360 179.360 ;
        RECT 99.380 177.660 99.520 182.780 ;
        RECT 104.380 182.500 104.640 182.760 ;
        RECT 103.520 182.440 104.640 182.500 ;
        RECT 103.520 182.360 104.580 182.440 ;
        RECT 99.780 179.380 100.040 179.700 ;
        RECT 102.080 179.380 102.340 179.700 ;
        RECT 99.840 178.340 99.980 179.380 ;
        RECT 99.780 178.020 100.040 178.340 ;
        RECT 102.140 177.660 102.280 179.380 ;
        RECT 98.400 177.340 98.660 177.660 ;
        RECT 99.320 177.340 99.580 177.660 ;
        RECT 102.080 177.340 102.340 177.660 ;
        RECT 91.800 175.785 93.680 176.155 ;
        RECT 98.460 174.600 98.600 177.340 ;
        RECT 100.700 176.320 100.960 176.640 ;
        RECT 102.080 176.320 102.340 176.640 ;
        RECT 98.400 174.280 98.660 174.600 ;
        RECT 98.460 173.920 98.600 174.280 ;
        RECT 98.400 173.600 98.660 173.920 ;
        RECT 91.040 172.580 91.300 172.900 ;
        RECT 98.400 171.560 98.660 171.880 ;
        RECT 89.660 170.880 89.920 171.200 ;
        RECT 89.720 169.840 89.860 170.880 ;
        RECT 91.800 170.345 93.680 170.715 ;
        RECT 98.460 170.180 98.600 171.560 ;
        RECT 98.400 169.860 98.660 170.180 ;
        RECT 89.660 169.520 89.920 169.840 ;
        RECT 91.960 169.180 92.220 169.500 ;
        RECT 87.820 168.840 88.080 169.160 ;
        RECT 91.040 168.840 91.300 169.160 ;
        RECT 84.140 168.500 84.400 168.820 ;
        RECT 84.200 167.120 84.340 168.500 ;
        RECT 84.140 166.800 84.400 167.120 ;
        RECT 83.740 166.040 84.340 166.180 ;
        RECT 83.220 163.400 83.480 163.720 ;
        RECT 80.980 160.660 81.120 162.720 ;
        RECT 81.900 162.640 83.880 162.780 ;
        RECT 82.760 161.700 83.020 162.020 ;
        RECT 80.920 160.340 81.180 160.660 ;
        RECT 80.980 159.300 81.120 160.340 ;
        RECT 80.920 158.980 81.180 159.300 ;
        RECT 81.370 159.125 81.650 159.495 ;
        RECT 80.980 156.240 81.120 158.980 ;
        RECT 80.920 155.920 81.180 156.240 ;
        RECT 80.520 155.160 81.120 155.300 ;
        RECT 80.460 154.560 80.720 154.880 ;
        RECT 80.000 150.140 80.260 150.460 ;
        RECT 79.540 149.800 79.800 150.120 ;
        RECT 78.160 149.460 78.420 149.780 ;
        RECT 78.220 148.080 78.360 149.460 ;
        RECT 80.060 148.420 80.200 150.140 ;
        RECT 80.000 148.100 80.260 148.420 ;
        RECT 78.160 147.760 78.420 148.080 ;
        RECT 78.160 147.080 78.420 147.400 ;
        RECT 80.000 147.080 80.260 147.400 ;
        RECT 78.220 146.720 78.360 147.080 ;
        RECT 78.160 146.400 78.420 146.720 ;
        RECT 79.540 146.400 79.800 146.720 ;
        RECT 76.800 145.865 78.680 146.235 ;
        RECT 79.600 145.360 79.740 146.400 ;
        RECT 79.540 145.040 79.800 145.360 ;
        RECT 76.800 140.425 78.680 140.795 ;
        RECT 80.060 139.920 80.200 147.080 ;
        RECT 80.000 139.600 80.260 139.920 ;
        RECT 79.540 138.240 79.800 138.560 ;
        RECT 79.600 136.520 79.740 138.240 ;
        RECT 80.000 137.220 80.260 137.540 ;
        RECT 76.320 136.200 76.580 136.520 ;
        RECT 79.540 136.200 79.800 136.520 ;
        RECT 79.080 135.520 79.340 135.840 ;
        RECT 76.800 134.985 78.680 135.355 ;
        RECT 79.140 134.480 79.280 135.520 ;
        RECT 79.080 134.160 79.340 134.480 ;
        RECT 80.060 132.100 80.200 137.220 ;
        RECT 80.520 134.140 80.660 154.560 ;
        RECT 80.980 145.700 81.120 155.160 ;
        RECT 80.920 145.380 81.180 145.700 ;
        RECT 81.440 145.020 81.580 159.125 ;
        RECT 81.840 157.960 82.100 158.280 ;
        RECT 81.900 155.900 82.040 157.960 ;
        RECT 82.300 157.620 82.560 157.940 ;
        RECT 82.360 155.900 82.500 157.620 ;
        RECT 82.820 155.900 82.960 161.700 ;
        RECT 83.220 160.000 83.480 160.320 ;
        RECT 83.280 157.940 83.420 160.000 ;
        RECT 83.220 157.620 83.480 157.940 ;
        RECT 81.840 155.580 82.100 155.900 ;
        RECT 82.300 155.580 82.560 155.900 ;
        RECT 82.760 155.580 83.020 155.900 ;
        RECT 82.360 155.220 82.500 155.580 ;
        RECT 82.300 154.900 82.560 155.220 ;
        RECT 81.840 149.120 82.100 149.440 ;
        RECT 81.380 144.700 81.640 145.020 ;
        RECT 80.920 143.680 81.180 144.000 ;
        RECT 80.460 133.820 80.720 134.140 ;
        RECT 80.980 133.540 81.120 143.680 ;
        RECT 81.380 139.940 81.640 140.260 ;
        RECT 81.440 136.520 81.580 139.940 ;
        RECT 81.380 136.200 81.640 136.520 ;
        RECT 80.520 133.400 81.120 133.540 ;
        RECT 80.000 131.780 80.260 132.100 ;
        RECT 80.000 130.760 80.260 131.080 ;
        RECT 76.800 129.545 78.680 129.915 ;
        RECT 78.620 128.040 78.880 128.360 ;
        RECT 78.680 126.660 78.820 128.040 ;
        RECT 79.080 127.700 79.340 128.020 ;
        RECT 79.140 126.660 79.280 127.700 ;
        RECT 78.620 126.340 78.880 126.660 ;
        RECT 79.080 126.340 79.340 126.660 ;
        RECT 76.800 124.105 78.680 124.475 ;
        RECT 79.140 119.520 79.280 126.340 ;
        RECT 79.540 125.660 79.800 125.980 ;
        RECT 79.600 120.540 79.740 125.660 ;
        RECT 79.540 120.220 79.800 120.540 ;
        RECT 79.540 119.770 79.800 119.860 ;
        RECT 80.060 119.770 80.200 130.760 ;
        RECT 80.520 129.040 80.660 133.400 ;
        RECT 80.460 128.720 80.720 129.040 ;
        RECT 80.460 128.040 80.720 128.360 ;
        RECT 80.520 126.660 80.660 128.040 ;
        RECT 81.900 127.680 82.040 149.120 ;
        RECT 83.220 147.760 83.480 148.080 ;
        RECT 83.280 147.400 83.420 147.760 ;
        RECT 82.300 147.080 82.560 147.400 ;
        RECT 83.220 147.080 83.480 147.400 ;
        RECT 82.360 146.720 82.500 147.080 ;
        RECT 82.760 146.740 83.020 147.060 ;
        RECT 82.300 146.400 82.560 146.720 ;
        RECT 82.300 139.150 82.560 139.240 ;
        RECT 82.820 139.150 82.960 146.740 ;
        RECT 83.280 139.240 83.420 147.080 ;
        RECT 82.300 139.010 82.960 139.150 ;
        RECT 82.300 138.920 82.560 139.010 ;
        RECT 83.220 138.920 83.480 139.240 ;
        RECT 82.360 137.200 82.500 138.920 ;
        RECT 82.300 136.880 82.560 137.200 ;
        RECT 83.280 136.520 83.420 138.920 ;
        RECT 83.220 136.200 83.480 136.520 ;
        RECT 83.740 133.800 83.880 162.640 ;
        RECT 84.200 136.180 84.340 166.040 ;
        RECT 87.880 164.740 88.020 168.840 ;
        RECT 88.740 166.460 89.000 166.780 ;
        RECT 87.820 164.420 88.080 164.740 ;
        RECT 88.800 160.660 88.940 166.460 ;
        RECT 91.100 166.440 91.240 168.840 ;
        RECT 92.020 166.440 92.160 169.180 ;
        RECT 100.240 166.800 100.500 167.120 ;
        RECT 91.040 166.120 91.300 166.440 ;
        RECT 91.960 166.120 92.220 166.440 ;
        RECT 93.800 166.120 94.060 166.440 ;
        RECT 94.720 166.120 94.980 166.440 ;
        RECT 98.400 166.120 98.660 166.440 ;
        RECT 91.100 163.040 91.240 166.120 ;
        RECT 92.020 165.760 92.160 166.120 ;
        RECT 91.960 165.440 92.220 165.760 ;
        RECT 91.800 164.905 93.680 165.275 ;
        RECT 93.860 164.060 94.000 166.120 ;
        RECT 93.800 163.740 94.060 164.060 ;
        RECT 91.040 162.720 91.300 163.040 ;
        RECT 88.740 160.340 89.000 160.660 ;
        RECT 88.280 160.000 88.540 160.320 ;
        RECT 84.590 158.445 84.870 158.815 ;
        RECT 88.340 158.620 88.480 160.000 ;
        RECT 88.800 158.620 88.940 160.340 ;
        RECT 84.660 155.900 84.800 158.445 ;
        RECT 88.280 158.300 88.540 158.620 ;
        RECT 88.740 158.300 89.000 158.620 ;
        RECT 91.100 158.280 91.240 162.720 ;
        RECT 94.780 162.020 94.920 166.120 ;
        RECT 96.560 165.440 96.820 165.760 ;
        RECT 94.720 161.700 94.980 162.020 ;
        RECT 94.260 161.360 94.520 161.680 ;
        RECT 91.800 159.465 93.680 159.835 ;
        RECT 94.320 159.300 94.460 161.360 ;
        RECT 94.260 158.980 94.520 159.300 ;
        RECT 96.620 158.280 96.760 165.440 ;
        RECT 98.460 163.380 98.600 166.120 ;
        RECT 98.400 163.060 98.660 163.380 ;
        RECT 97.480 162.720 97.740 163.040 ;
        RECT 97.540 161.340 97.680 162.720 ;
        RECT 97.480 161.020 97.740 161.340 ;
        RECT 97.020 160.680 97.280 161.000 ;
        RECT 97.080 159.300 97.220 160.680 ;
        RECT 97.020 158.980 97.280 159.300 ;
        RECT 91.040 157.960 91.300 158.280 ;
        RECT 96.560 157.960 96.820 158.280 ;
        RECT 84.600 155.580 84.860 155.900 ;
        RECT 91.100 153.770 91.240 157.960 ;
        RECT 95.180 157.620 95.440 157.940 ;
        RECT 91.800 154.025 93.680 154.395 ;
        RECT 91.100 153.630 92.160 153.770 ;
        RECT 92.020 153.180 92.160 153.630 ;
        RECT 91.960 152.860 92.220 153.180 ;
        RECT 93.800 153.090 94.060 153.180 ;
        RECT 93.400 152.950 94.060 153.090 ;
        RECT 87.820 152.180 88.080 152.500 ;
        RECT 86.440 151.840 86.700 152.160 ;
        RECT 86.500 151.140 86.640 151.840 ;
        RECT 86.440 150.820 86.700 151.140 ;
        RECT 85.980 150.140 86.240 150.460 ;
        RECT 85.060 149.800 85.320 150.120 ;
        RECT 85.120 148.420 85.260 149.800 ;
        RECT 85.060 148.100 85.320 148.420 ;
        RECT 84.600 144.700 84.860 145.020 ;
        RECT 84.660 140.260 84.800 144.700 ;
        RECT 85.120 144.680 85.260 148.100 ;
        RECT 86.040 146.720 86.180 150.140 ;
        RECT 86.500 147.740 86.640 150.820 ;
        RECT 87.880 150.655 88.020 152.180 ;
        RECT 93.400 151.140 93.540 152.950 ;
        RECT 93.800 152.860 94.060 152.950 ;
        RECT 93.800 151.840 94.060 152.160 ;
        RECT 93.860 151.140 94.000 151.840 ;
        RECT 93.340 150.820 93.600 151.140 ;
        RECT 93.800 150.820 94.060 151.140 ;
        RECT 87.810 150.285 88.090 150.655 ;
        RECT 93.800 149.460 94.060 149.780 ;
        RECT 94.260 149.460 94.520 149.780 ;
        RECT 90.580 149.120 90.840 149.440 ;
        RECT 86.440 147.420 86.700 147.740 ;
        RECT 90.640 147.060 90.780 149.120 ;
        RECT 91.800 148.585 93.680 148.955 ;
        RECT 91.040 147.420 91.300 147.740 ;
        RECT 90.580 146.740 90.840 147.060 ;
        RECT 85.980 146.400 86.240 146.720 ;
        RECT 86.040 145.700 86.180 146.400 ;
        RECT 91.100 145.700 91.240 147.420 ;
        RECT 93.860 147.060 94.000 149.460 ;
        RECT 94.320 147.400 94.460 149.460 ;
        RECT 95.240 147.400 95.380 157.620 ;
        RECT 98.460 155.900 98.600 163.060 ;
        RECT 100.300 159.300 100.440 166.800 ;
        RECT 100.240 158.980 100.500 159.300 ;
        RECT 98.400 155.580 98.660 155.900 ;
        RECT 98.860 155.580 99.120 155.900 ;
        RECT 98.920 153.860 99.060 155.580 ;
        RECT 99.780 154.560 100.040 154.880 ;
        RECT 98.860 153.540 99.120 153.860 ;
        RECT 95.640 150.480 95.900 150.800 ;
        RECT 95.700 148.420 95.840 150.480 ;
        RECT 99.310 150.285 99.590 150.655 ;
        RECT 96.560 149.120 96.820 149.440 ;
        RECT 96.620 148.420 96.760 149.120 ;
        RECT 95.640 148.100 95.900 148.420 ;
        RECT 96.560 148.100 96.820 148.420 ;
        RECT 94.260 147.080 94.520 147.400 ;
        RECT 95.180 147.080 95.440 147.400 ;
        RECT 93.800 146.740 94.060 147.060 ;
        RECT 85.980 145.380 86.240 145.700 ;
        RECT 91.040 145.380 91.300 145.700 ;
        RECT 85.060 144.360 85.320 144.680 ;
        RECT 84.600 139.940 84.860 140.260 ;
        RECT 84.660 137.540 84.800 139.940 ;
        RECT 85.120 139.240 85.260 144.360 ;
        RECT 91.800 143.145 93.680 143.515 ;
        RECT 86.440 139.260 86.700 139.580 ;
        RECT 85.060 138.920 85.320 139.240 ;
        RECT 85.120 137.540 85.260 138.920 ;
        RECT 84.600 137.220 84.860 137.540 ;
        RECT 85.060 137.220 85.320 137.540 ;
        RECT 86.500 136.860 86.640 139.260 ;
        RECT 94.320 138.900 94.460 147.080 ;
        RECT 96.620 145.020 96.760 148.100 ;
        RECT 97.020 146.400 97.280 146.720 ;
        RECT 97.080 145.700 97.220 146.400 ;
        RECT 97.020 145.380 97.280 145.700 ;
        RECT 96.560 144.700 96.820 145.020 ;
        RECT 98.860 138.920 99.120 139.240 ;
        RECT 94.260 138.580 94.520 138.900 ;
        RECT 91.040 138.240 91.300 138.560 ;
        RECT 86.900 136.880 87.160 137.200 ;
        RECT 86.440 136.540 86.700 136.860 ;
        RECT 84.140 135.860 84.400 136.180 ;
        RECT 85.060 135.520 85.320 135.840 ;
        RECT 85.120 134.480 85.260 135.520 ;
        RECT 85.060 134.160 85.320 134.480 ;
        RECT 86.500 133.800 86.640 136.540 ;
        RECT 83.680 133.480 83.940 133.800 ;
        RECT 86.440 133.480 86.700 133.800 ;
        RECT 83.220 132.800 83.480 133.120 ;
        RECT 83.280 129.380 83.420 132.800 ;
        RECT 83.220 129.060 83.480 129.380 ;
        RECT 81.840 127.360 82.100 127.680 ;
        RECT 83.680 127.360 83.940 127.680 ;
        RECT 84.600 127.360 84.860 127.680 ;
        RECT 80.460 126.340 80.720 126.660 ;
        RECT 82.760 124.980 83.020 125.300 ;
        RECT 82.820 123.940 82.960 124.980 ;
        RECT 82.760 123.620 83.020 123.940 ;
        RECT 83.740 123.260 83.880 127.360 ;
        RECT 84.660 125.980 84.800 127.360 ;
        RECT 84.600 125.660 84.860 125.980 ;
        RECT 85.520 125.320 85.780 125.640 ;
        RECT 85.580 123.940 85.720 125.320 ;
        RECT 85.520 123.620 85.780 123.940 ;
        RECT 83.220 122.940 83.480 123.260 ;
        RECT 83.680 122.940 83.940 123.260 ;
        RECT 83.280 120.200 83.420 122.940 ;
        RECT 83.680 120.220 83.940 120.540 ;
        RECT 83.220 119.880 83.480 120.200 ;
        RECT 79.540 119.630 80.200 119.770 ;
        RECT 79.540 119.540 79.800 119.630 ;
        RECT 79.080 119.200 79.340 119.520 ;
        RECT 76.800 118.665 78.680 119.035 ;
        RECT 79.140 118.500 79.280 119.200 ;
        RECT 79.080 118.180 79.340 118.500 ;
        RECT 79.600 117.480 79.740 119.540 ;
        RECT 80.920 119.200 81.180 119.520 ;
        RECT 82.760 119.200 83.020 119.520 ;
        RECT 80.980 117.820 81.120 119.200 ;
        RECT 80.920 117.500 81.180 117.820 ;
        RECT 79.540 117.160 79.800 117.480 ;
        RECT 79.600 115.780 79.740 117.160 ;
        RECT 79.540 115.460 79.800 115.780 ;
        RECT 82.820 114.420 82.960 119.200 ;
        RECT 83.280 118.160 83.420 119.880 ;
        RECT 83.220 117.840 83.480 118.160 ;
        RECT 83.740 117.140 83.880 120.220 ;
        RECT 84.140 119.880 84.400 120.200 ;
        RECT 84.200 118.500 84.340 119.880 ;
        RECT 84.600 119.200 84.860 119.520 ;
        RECT 84.140 118.180 84.400 118.500 ;
        RECT 83.680 116.820 83.940 117.140 ;
        RECT 84.660 115.100 84.800 119.200 ;
        RECT 85.520 117.160 85.780 117.480 ;
        RECT 85.580 115.100 85.720 117.160 ;
        RECT 84.600 114.780 84.860 115.100 ;
        RECT 85.520 114.780 85.780 115.100 ;
        RECT 86.440 114.780 86.700 115.100 ;
        RECT 82.760 114.100 83.020 114.420 ;
        RECT 76.800 113.225 78.680 113.595 ;
        RECT 78.160 112.060 78.420 112.380 ;
        RECT 81.380 112.060 81.640 112.380 ;
        RECT 78.220 109.320 78.360 112.060 ;
        RECT 81.440 109.660 81.580 112.060 ;
        RECT 81.840 111.720 82.100 112.040 ;
        RECT 81.380 109.340 81.640 109.660 ;
        RECT 78.160 109.000 78.420 109.320 ;
        RECT 79.080 109.000 79.340 109.320 ;
        RECT 75.860 108.660 76.120 108.980 ;
        RECT 76.800 107.785 78.680 108.155 ;
        RECT 74.940 106.620 75.200 106.940 ;
        RECT 68.500 106.510 68.760 106.600 ;
        RECT 68.100 106.370 68.760 106.510 ;
        RECT 64.360 105.940 64.620 106.260 ;
        RECT 63.900 105.600 64.160 105.920 ;
        RECT 61.800 105.065 63.680 105.435 ;
        RECT 63.960 104.220 64.100 105.600 ;
        RECT 52.400 103.560 52.660 103.880 ;
        RECT 56.600 103.540 56.740 104.160 ;
        RECT 57.920 103.900 58.180 104.220 ;
        RECT 63.900 103.900 64.160 104.220 ;
        RECT 64.420 103.540 64.560 105.940 ;
        RECT 54.700 103.220 54.960 103.540 ;
        RECT 56.540 103.220 56.800 103.540 ;
        RECT 61.140 103.220 61.400 103.540 ;
        RECT 64.360 103.220 64.620 103.540 ;
        RECT 50.090 89.040 50.370 89.210 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 54.760 88.660 54.900 103.220 ;
        RECT 61.200 98.860 61.340 103.220 ;
        RECT 61.800 99.625 63.680 99.995 ;
        RECT 61.200 98.720 62.260 98.860 ;
        RECT 62.120 89.210 62.260 98.720 ;
        RECT 68.100 89.840 68.240 106.370 ;
        RECT 68.500 106.280 68.760 106.370 ;
        RECT 73.560 106.280 73.820 106.600 ;
        RECT 73.620 104.900 73.760 106.280 ;
        RECT 75.860 105.600 76.120 105.920 ;
        RECT 73.560 104.580 73.820 104.900 ;
        RECT 73.620 104.220 73.760 104.580 ;
        RECT 75.920 104.220 76.060 105.600 ;
        RECT 79.140 104.900 79.280 109.000 ;
        RECT 79.540 108.320 79.800 108.640 ;
        RECT 79.080 104.580 79.340 104.900 ;
        RECT 73.560 103.900 73.820 104.220 ;
        RECT 75.860 103.900 76.120 104.220 ;
        RECT 79.600 103.880 79.740 108.320 ;
        RECT 81.900 107.280 82.040 111.720 ;
        RECT 83.680 108.320 83.940 108.640 ;
        RECT 83.740 107.280 83.880 108.320 ;
        RECT 81.840 106.960 82.100 107.280 ;
        RECT 83.680 106.960 83.940 107.280 ;
        RECT 86.500 106.600 86.640 114.780 ;
        RECT 86.960 106.940 87.100 136.880 ;
        RECT 91.100 136.860 91.240 138.240 ;
        RECT 91.800 137.705 93.680 138.075 ;
        RECT 91.040 136.540 91.300 136.860 ;
        RECT 91.500 136.540 91.760 136.860 ;
        RECT 88.280 135.860 88.540 136.180 ;
        RECT 88.340 134.820 88.480 135.860 ;
        RECT 88.280 134.500 88.540 134.820 ;
        RECT 90.580 134.160 90.840 134.480 ;
        RECT 88.280 133.820 88.540 134.140 ;
        RECT 88.340 131.080 88.480 133.820 ;
        RECT 90.640 132.100 90.780 134.160 ;
        RECT 91.560 133.800 91.700 136.540 ;
        RECT 93.340 136.430 93.600 136.520 ;
        RECT 92.940 136.290 93.600 136.430 ;
        RECT 92.940 135.840 93.080 136.290 ;
        RECT 93.340 136.200 93.600 136.290 ;
        RECT 94.320 136.180 94.460 138.580 ;
        RECT 98.400 138.240 98.660 138.560 ;
        RECT 97.940 136.200 98.200 136.520 ;
        RECT 94.260 135.860 94.520 136.180 ;
        RECT 92.880 135.520 93.140 135.840 ;
        RECT 93.800 135.520 94.060 135.840 ;
        RECT 91.500 133.480 91.760 133.800 ;
        RECT 91.800 132.265 93.680 132.635 ;
        RECT 90.580 131.780 90.840 132.100 ;
        RECT 88.280 130.760 88.540 131.080 ;
        RECT 91.040 130.760 91.300 131.080 ;
        RECT 88.280 129.060 88.540 129.380 ;
        RECT 88.340 125.980 88.480 129.060 ;
        RECT 88.280 125.660 88.540 125.980 ;
        RECT 91.100 123.260 91.240 130.760 ;
        RECT 93.860 128.700 94.000 135.520 ;
        RECT 98.000 134.140 98.140 136.200 ;
        RECT 98.460 136.180 98.600 138.240 ;
        RECT 98.920 136.520 99.060 138.920 ;
        RECT 99.380 136.520 99.520 150.285 ;
        RECT 98.860 136.200 99.120 136.520 ;
        RECT 99.320 136.200 99.580 136.520 ;
        RECT 98.400 135.860 98.660 136.180 ;
        RECT 98.460 134.140 98.600 135.860 ;
        RECT 99.380 134.335 99.520 136.200 ;
        RECT 97.940 133.820 98.200 134.140 ;
        RECT 98.400 133.820 98.660 134.140 ;
        RECT 99.310 133.965 99.590 134.335 ;
        RECT 99.840 134.140 99.980 154.560 ;
        RECT 100.240 136.200 100.500 136.520 ;
        RECT 100.300 134.820 100.440 136.200 ;
        RECT 100.240 134.500 100.500 134.820 ;
        RECT 99.780 133.820 100.040 134.140 ;
        RECT 95.180 133.480 95.440 133.800 ;
        RECT 94.720 132.800 94.980 133.120 ;
        RECT 93.800 128.380 94.060 128.700 ;
        RECT 91.560 128.020 94.000 128.100 ;
        RECT 91.500 127.960 94.000 128.020 ;
        RECT 91.500 127.700 91.760 127.960 ;
        RECT 91.800 126.825 93.680 127.195 ;
        RECT 93.340 124.980 93.600 125.300 ;
        RECT 93.400 123.940 93.540 124.980 ;
        RECT 93.340 123.620 93.600 123.940 ;
        RECT 91.040 122.940 91.300 123.260 ;
        RECT 91.800 121.385 93.680 121.755 ;
        RECT 93.340 119.880 93.600 120.200 ;
        RECT 87.360 119.200 87.620 119.520 ;
        RECT 87.420 117.820 87.560 119.200 ;
        RECT 93.400 118.500 93.540 119.880 ;
        RECT 93.860 119.520 94.000 127.960 ;
        RECT 93.800 119.200 94.060 119.520 ;
        RECT 93.340 118.180 93.600 118.500 ;
        RECT 87.360 117.500 87.620 117.820 ;
        RECT 93.860 117.480 94.000 119.200 ;
        RECT 93.800 117.160 94.060 117.480 ;
        RECT 88.280 116.480 88.540 116.800 ;
        RECT 91.040 116.480 91.300 116.800 ;
        RECT 88.340 115.100 88.480 116.480 ;
        RECT 88.280 114.780 88.540 115.100 ;
        RECT 91.100 114.420 91.240 116.480 ;
        RECT 91.800 115.945 93.680 116.315 ;
        RECT 93.860 115.780 94.000 117.160 ;
        RECT 93.800 115.460 94.060 115.780 ;
        RECT 91.040 114.100 91.300 114.420 ;
        RECT 92.870 112.885 93.150 113.255 ;
        RECT 92.940 112.720 93.080 112.885 ;
        RECT 92.880 112.400 93.140 112.720 ;
        RECT 91.800 110.505 93.680 110.875 ;
        RECT 94.780 109.320 94.920 132.800 ;
        RECT 95.240 129.380 95.380 133.480 ;
        RECT 98.460 131.080 98.600 133.820 ;
        RECT 100.760 133.800 100.900 176.320 ;
        RECT 101.150 163.885 101.430 164.255 ;
        RECT 101.220 163.720 101.360 163.885 ;
        RECT 101.160 163.400 101.420 163.720 ;
        RECT 101.620 151.840 101.880 152.160 ;
        RECT 101.160 135.520 101.420 135.840 ;
        RECT 101.220 134.480 101.360 135.520 ;
        RECT 101.160 134.160 101.420 134.480 ;
        RECT 100.700 133.480 100.960 133.800 ;
        RECT 99.780 132.800 100.040 133.120 ;
        RECT 101.160 132.800 101.420 133.120 ;
        RECT 98.400 130.760 98.660 131.080 ;
        RECT 95.180 129.060 95.440 129.380 ;
        RECT 95.630 129.205 95.910 129.575 ;
        RECT 98.460 129.380 98.600 130.760 ;
        RECT 95.700 129.040 95.840 129.205 ;
        RECT 98.400 129.060 98.660 129.380 ;
        RECT 95.640 128.720 95.900 129.040 ;
        RECT 98.460 125.980 98.600 129.060 ;
        RECT 98.860 128.040 99.120 128.360 ;
        RECT 98.920 126.660 99.060 128.040 ;
        RECT 98.860 126.340 99.120 126.660 ;
        RECT 98.400 125.660 98.660 125.980 ;
        RECT 99.320 125.320 99.580 125.640 ;
        RECT 99.380 120.200 99.520 125.320 ;
        RECT 99.320 119.880 99.580 120.200 ;
        RECT 99.840 109.320 99.980 132.800 ;
        RECT 100.240 131.440 100.500 131.760 ;
        RECT 100.300 128.700 100.440 131.440 ;
        RECT 100.240 128.380 100.500 128.700 ;
        RECT 100.300 125.640 100.440 128.380 ;
        RECT 101.220 125.640 101.360 132.800 ;
        RECT 100.240 125.320 100.500 125.640 ;
        RECT 101.160 125.320 101.420 125.640 ;
        RECT 100.240 122.940 100.500 123.260 ;
        RECT 100.300 120.200 100.440 122.940 ;
        RECT 100.240 119.880 100.500 120.200 ;
        RECT 101.160 119.200 101.420 119.520 ;
        RECT 100.240 117.160 100.500 117.480 ;
        RECT 100.300 115.780 100.440 117.160 ;
        RECT 100.240 115.460 100.500 115.780 ;
        RECT 101.220 114.760 101.360 119.200 ;
        RECT 101.160 114.440 101.420 114.760 ;
        RECT 101.680 114.080 101.820 151.840 ;
        RECT 102.140 133.800 102.280 176.320 ;
        RECT 102.540 168.160 102.800 168.480 ;
        RECT 102.600 161.340 102.740 168.160 ;
        RECT 102.540 161.020 102.800 161.340 ;
        RECT 102.600 160.180 102.740 161.020 ;
        RECT 102.600 160.040 103.200 160.180 ;
        RECT 102.540 156.260 102.800 156.580 ;
        RECT 102.600 155.220 102.740 156.260 ;
        RECT 103.060 156.240 103.200 160.040 ;
        RECT 103.000 155.920 103.260 156.240 ;
        RECT 102.540 154.900 102.800 155.220 ;
        RECT 103.000 153.770 103.260 153.860 ;
        RECT 102.600 153.630 103.260 153.770 ;
        RECT 102.600 147.140 102.740 153.630 ;
        RECT 103.000 153.540 103.260 153.630 ;
        RECT 103.520 151.220 103.660 182.360 ;
        RECT 104.840 181.760 105.100 182.080 ;
        RECT 104.900 180.380 105.040 181.760 ;
        RECT 104.840 180.060 105.100 180.380 ;
        RECT 104.840 174.510 105.100 174.600 ;
        RECT 105.360 174.510 105.500 185.500 ;
        RECT 105.760 185.160 106.020 185.480 ;
        RECT 105.820 183.780 105.960 185.160 ;
        RECT 106.800 183.945 108.680 184.315 ;
        RECT 105.760 183.460 106.020 183.780 ;
        RECT 105.760 182.780 106.020 183.100 ;
        RECT 106.220 182.780 106.480 183.100 ;
        RECT 108.060 182.780 108.320 183.100 ;
        RECT 109.440 182.780 109.700 183.100 ;
        RECT 105.820 181.060 105.960 182.780 ;
        RECT 105.760 180.740 106.020 181.060 ;
        RECT 105.760 180.060 106.020 180.380 ;
        RECT 105.820 177.320 105.960 180.060 ;
        RECT 106.280 177.570 106.420 182.780 ;
        RECT 108.120 180.380 108.260 182.780 ;
        RECT 108.060 180.060 108.320 180.380 ;
        RECT 108.980 179.720 109.240 180.040 ;
        RECT 106.800 178.505 108.680 178.875 ;
        RECT 109.040 178.000 109.180 179.720 ;
        RECT 108.980 177.680 109.240 178.000 ;
        RECT 109.500 177.660 109.640 182.780 ;
        RECT 106.680 177.570 106.940 177.660 ;
        RECT 106.280 177.430 106.940 177.570 ;
        RECT 106.680 177.340 106.940 177.430 ;
        RECT 108.060 177.340 108.320 177.660 ;
        RECT 109.440 177.340 109.700 177.660 ;
        RECT 105.760 177.000 106.020 177.320 ;
        RECT 105.820 174.600 105.960 177.000 ;
        RECT 106.220 175.300 106.480 175.620 ;
        RECT 104.840 174.370 105.500 174.510 ;
        RECT 104.840 174.280 105.100 174.370 ;
        RECT 105.760 174.280 106.020 174.600 ;
        RECT 104.380 173.940 104.640 174.260 ;
        RECT 103.920 154.560 104.180 154.880 ;
        RECT 103.060 151.080 103.660 151.220 ;
        RECT 103.060 147.740 103.200 151.080 ;
        RECT 103.460 150.480 103.720 150.800 ;
        RECT 103.520 148.420 103.660 150.480 ;
        RECT 103.460 148.100 103.720 148.420 ;
        RECT 103.000 147.420 103.260 147.740 ;
        RECT 102.600 147.000 103.200 147.140 ;
        RECT 102.540 139.600 102.800 139.920 ;
        RECT 102.600 134.820 102.740 139.600 ;
        RECT 102.540 134.500 102.800 134.820 ;
        RECT 102.540 133.820 102.800 134.140 ;
        RECT 102.080 133.480 102.340 133.800 ;
        RECT 102.600 131.760 102.740 133.820 ;
        RECT 102.540 131.440 102.800 131.760 ;
        RECT 103.060 128.020 103.200 147.000 ;
        RECT 103.980 134.140 104.120 154.560 ;
        RECT 104.440 153.180 104.580 173.940 ;
        RECT 106.280 172.560 106.420 175.300 ;
        RECT 106.740 174.940 106.880 177.340 ;
        RECT 108.120 175.620 108.260 177.340 ;
        RECT 108.060 175.300 108.320 175.620 ;
        RECT 108.980 174.960 109.240 175.280 ;
        RECT 106.680 174.620 106.940 174.940 ;
        RECT 106.800 173.065 108.680 173.435 ;
        RECT 106.220 172.240 106.480 172.560 ;
        RECT 105.760 171.560 106.020 171.880 ;
        RECT 105.820 166.440 105.960 171.560 ;
        RECT 107.140 170.880 107.400 171.200 ;
        RECT 107.200 168.820 107.340 170.880 ;
        RECT 107.140 168.500 107.400 168.820 ;
        RECT 106.800 167.625 108.680 167.995 ;
        RECT 104.840 166.120 105.100 166.440 ;
        RECT 105.760 166.120 106.020 166.440 ;
        RECT 104.900 159.300 105.040 166.120 ;
        RECT 105.300 162.720 105.560 163.040 ;
        RECT 104.840 158.980 105.100 159.300 ;
        RECT 105.360 158.280 105.500 162.720 ;
        RECT 105.820 161.000 105.960 166.120 ;
        RECT 109.040 166.100 109.180 174.960 ;
        RECT 109.960 174.600 110.100 188.220 ;
        RECT 110.360 185.160 110.620 185.480 ;
        RECT 110.420 182.420 110.560 185.160 ;
        RECT 110.880 182.760 111.020 193.320 ;
        RECT 112.200 192.980 112.460 193.300 ;
        RECT 112.260 185.140 112.400 192.980 ;
        RECT 112.720 191.940 112.860 194.340 ;
        RECT 115.880 193.660 116.140 193.980 ;
        RECT 112.660 191.620 112.920 191.940 ;
        RECT 113.120 189.920 113.380 190.240 ;
        RECT 113.180 188.540 113.320 189.920 ;
        RECT 113.120 188.220 113.380 188.540 ;
        RECT 112.200 184.820 112.460 185.140 ;
        RECT 111.740 184.480 112.000 184.800 ;
        RECT 111.800 183.100 111.940 184.480 ;
        RECT 111.740 182.780 112.000 183.100 ;
        RECT 110.820 182.440 111.080 182.760 ;
        RECT 110.360 182.100 110.620 182.420 ;
        RECT 109.440 174.280 109.700 174.600 ;
        RECT 109.900 174.280 110.160 174.600 ;
        RECT 109.500 172.220 109.640 174.280 ;
        RECT 109.900 173.600 110.160 173.920 ;
        RECT 109.960 172.220 110.100 173.600 ;
        RECT 110.420 172.560 110.560 182.100 ;
        RECT 110.880 177.320 111.020 182.440 ;
        RECT 111.800 178.340 111.940 182.780 ;
        RECT 112.260 178.340 112.400 184.820 ;
        RECT 115.940 180.380 116.080 193.660 ;
        RECT 117.780 191.940 117.920 195.700 ;
        RECT 118.240 194.320 118.380 195.700 ;
        RECT 118.180 194.000 118.440 194.320 ;
        RECT 117.720 191.620 117.980 191.940 ;
        RECT 118.240 190.920 118.380 194.000 ;
        RECT 119.100 192.640 119.360 192.960 ;
        RECT 119.160 190.920 119.300 192.640 ;
        RECT 121.800 192.105 123.680 192.475 ;
        RECT 118.180 190.600 118.440 190.920 ;
        RECT 119.100 190.600 119.360 190.920 ;
        RECT 116.340 190.260 116.600 190.580 ;
        RECT 116.400 189.220 116.540 190.260 ;
        RECT 116.340 188.900 116.600 189.220 ;
        RECT 118.240 188.200 118.380 190.600 ;
        RECT 118.180 187.880 118.440 188.200 ;
        RECT 117.720 182.780 117.980 183.100 ;
        RECT 116.800 181.760 117.060 182.080 ;
        RECT 115.880 180.060 116.140 180.380 ;
        RECT 111.740 178.020 112.000 178.340 ;
        RECT 112.200 178.020 112.460 178.340 ;
        RECT 116.860 177.660 117.000 181.760 ;
        RECT 117.780 181.060 117.920 182.780 ;
        RECT 118.240 182.760 118.380 187.880 ;
        RECT 121.800 186.665 123.680 187.035 ;
        RECT 124.620 183.120 124.880 183.440 ;
        RECT 118.180 182.440 118.440 182.760 ;
        RECT 117.720 180.740 117.980 181.060 ;
        RECT 118.240 179.360 118.380 182.440 ;
        RECT 121.800 181.225 123.680 181.595 ;
        RECT 124.680 181.060 124.820 183.120 ;
        RECT 124.620 180.740 124.880 181.060 ;
        RECT 121.860 179.720 122.120 180.040 ;
        RECT 118.640 179.380 118.900 179.700 ;
        RECT 118.180 179.040 118.440 179.360 ;
        RECT 118.700 178.340 118.840 179.380 ;
        RECT 118.640 178.020 118.900 178.340 ;
        RECT 121.920 178.000 122.060 179.720 ;
        RECT 121.860 177.680 122.120 178.000 ;
        RECT 116.800 177.340 117.060 177.660 ;
        RECT 110.820 177.000 111.080 177.320 ;
        RECT 121.800 175.785 123.680 176.155 ;
        RECT 119.100 174.280 119.360 174.600 ;
        RECT 118.180 173.600 118.440 173.920 ;
        RECT 118.240 172.560 118.380 173.600 ;
        RECT 119.160 172.900 119.300 174.280 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 119.100 172.580 119.360 172.900 ;
        RECT 110.360 172.240 110.620 172.560 ;
        RECT 118.180 172.240 118.440 172.560 ;
        RECT 109.440 171.900 109.700 172.220 ;
        RECT 109.900 171.900 110.160 172.220 ;
        RECT 114.500 171.220 114.760 171.540 ;
        RECT 111.280 170.880 111.540 171.200 ;
        RECT 113.580 170.880 113.840 171.200 ;
        RECT 109.900 169.180 110.160 169.500 ;
        RECT 108.980 165.780 109.240 166.100 ;
        RECT 109.960 164.820 110.100 169.180 ;
        RECT 110.360 168.500 110.620 168.820 ;
        RECT 110.420 167.460 110.560 168.500 ;
        RECT 110.820 168.160 111.080 168.480 ;
        RECT 110.360 167.140 110.620 167.460 ;
        RECT 110.880 166.780 111.020 168.160 ;
        RECT 110.820 166.460 111.080 166.780 ;
        RECT 110.820 165.780 111.080 166.100 ;
        RECT 109.500 164.680 110.100 164.820 ;
        RECT 108.980 164.080 109.240 164.400 ;
        RECT 106.220 163.060 106.480 163.380 ;
        RECT 106.280 162.020 106.420 163.060 ;
        RECT 106.800 162.185 108.680 162.555 ;
        RECT 106.220 161.700 106.480 162.020 ;
        RECT 105.760 160.680 106.020 161.000 ;
        RECT 109.040 158.280 109.180 164.080 ;
        RECT 109.500 158.960 109.640 164.680 ;
        RECT 110.360 163.740 110.620 164.060 ;
        RECT 109.900 162.720 110.160 163.040 ;
        RECT 109.960 162.020 110.100 162.720 ;
        RECT 109.900 161.700 110.160 162.020 ;
        RECT 110.420 161.340 110.560 163.740 ;
        RECT 110.360 161.020 110.620 161.340 ;
        RECT 110.880 160.740 111.020 165.780 ;
        RECT 110.420 160.600 111.020 160.740 ;
        RECT 109.440 158.640 109.700 158.960 ;
        RECT 105.300 157.960 105.560 158.280 ;
        RECT 108.980 157.960 109.240 158.280 ;
        RECT 109.440 157.960 109.700 158.280 ;
        RECT 109.900 157.960 110.160 158.280 ;
        RECT 108.980 157.280 109.240 157.600 ;
        RECT 106.800 156.745 108.680 157.115 ;
        RECT 108.520 156.260 108.780 156.580 ;
        RECT 105.300 155.580 105.560 155.900 ;
        RECT 105.360 153.520 105.500 155.580 ;
        RECT 106.680 154.560 106.940 154.880 ;
        RECT 105.300 153.200 105.560 153.520 ;
        RECT 104.380 152.860 104.640 153.180 ;
        RECT 106.740 152.840 106.880 154.560 ;
        RECT 108.060 153.200 108.320 153.520 ;
        RECT 106.680 152.520 106.940 152.840 ;
        RECT 107.600 152.750 107.860 152.840 ;
        RECT 108.120 152.750 108.260 153.200 ;
        RECT 108.580 152.840 108.720 156.260 ;
        RECT 107.600 152.610 108.260 152.750 ;
        RECT 107.600 152.520 107.860 152.610 ;
        RECT 108.520 152.520 108.780 152.840 ;
        RECT 104.840 152.180 105.100 152.500 ;
        RECT 104.900 151.140 105.040 152.180 ;
        RECT 108.580 152.160 108.720 152.520 ;
        RECT 105.300 151.840 105.560 152.160 ;
        RECT 108.520 151.840 108.780 152.160 ;
        RECT 104.840 150.820 105.100 151.140 ;
        RECT 104.380 148.100 104.640 148.420 ;
        RECT 103.920 133.820 104.180 134.140 ;
        RECT 103.460 132.800 103.720 133.120 ;
        RECT 103.000 127.700 103.260 128.020 ;
        RECT 102.540 119.540 102.800 119.860 ;
        RECT 102.600 118.500 102.740 119.540 ;
        RECT 102.540 118.180 102.800 118.500 ;
        RECT 101.620 113.760 101.880 114.080 ;
        RECT 103.520 109.320 103.660 132.800 ;
        RECT 104.440 112.040 104.580 148.100 ;
        RECT 105.360 147.400 105.500 151.840 ;
        RECT 106.800 151.305 108.680 151.675 ;
        RECT 107.590 150.285 107.870 150.655 ;
        RECT 107.660 150.120 107.800 150.285 ;
        RECT 108.060 150.140 108.320 150.460 ;
        RECT 107.600 149.800 107.860 150.120 ;
        RECT 106.220 148.100 106.480 148.420 ;
        RECT 105.300 147.080 105.560 147.400 ;
        RECT 105.300 138.920 105.560 139.240 ;
        RECT 105.360 137.540 105.500 138.920 ;
        RECT 105.300 137.220 105.560 137.540 ;
        RECT 104.840 132.800 105.100 133.120 ;
        RECT 104.900 129.380 105.040 132.800 ;
        RECT 106.280 129.380 106.420 148.100 ;
        RECT 107.660 147.740 107.800 149.800 ;
        RECT 107.600 147.420 107.860 147.740 ;
        RECT 108.120 147.400 108.260 150.140 ;
        RECT 108.060 147.080 108.320 147.400 ;
        RECT 108.120 146.720 108.260 147.080 ;
        RECT 108.060 146.400 108.320 146.720 ;
        RECT 106.800 145.865 108.680 146.235 ;
        RECT 109.040 145.020 109.180 157.280 ;
        RECT 109.500 155.900 109.640 157.960 ;
        RECT 109.440 155.580 109.700 155.900 ;
        RECT 109.500 152.840 109.640 155.580 ;
        RECT 109.960 153.860 110.100 157.960 ;
        RECT 109.900 153.540 110.160 153.860 ;
        RECT 109.960 153.180 110.100 153.540 ;
        RECT 109.900 152.860 110.160 153.180 ;
        RECT 109.440 152.520 109.700 152.840 ;
        RECT 109.900 150.140 110.160 150.460 ;
        RECT 109.960 147.400 110.100 150.140 ;
        RECT 109.900 147.080 110.160 147.400 ;
        RECT 109.440 146.400 109.700 146.720 ;
        RECT 109.500 145.020 109.640 146.400 ;
        RECT 108.980 144.700 109.240 145.020 ;
        RECT 109.440 144.700 109.700 145.020 ;
        RECT 109.960 144.420 110.100 147.080 ;
        RECT 110.420 144.680 110.560 160.600 ;
        RECT 110.820 160.000 111.080 160.320 ;
        RECT 110.880 156.240 111.020 160.000 ;
        RECT 110.820 155.920 111.080 156.240 ;
        RECT 110.820 154.560 111.080 154.880 ;
        RECT 108.980 144.020 109.240 144.340 ;
        RECT 109.500 144.280 110.100 144.420 ;
        RECT 110.360 144.360 110.620 144.680 ;
        RECT 109.040 142.980 109.180 144.020 ;
        RECT 108.980 142.660 109.240 142.980 ;
        RECT 106.800 140.425 108.680 140.795 ;
        RECT 109.500 139.580 109.640 144.280 ;
        RECT 109.900 143.680 110.160 144.000 ;
        RECT 110.360 143.680 110.620 144.000 ;
        RECT 109.440 139.260 109.700 139.580 ;
        RECT 108.980 135.860 109.240 136.180 ;
        RECT 106.800 134.985 108.680 135.355 ;
        RECT 108.050 133.965 108.330 134.335 ;
        RECT 109.040 134.140 109.180 135.860 ;
        RECT 109.500 134.140 109.640 139.260 ;
        RECT 108.060 133.820 108.320 133.965 ;
        RECT 108.980 133.820 109.240 134.140 ;
        RECT 109.440 133.820 109.700 134.140 ;
        RECT 109.960 132.100 110.100 143.680 ;
        RECT 110.420 139.920 110.560 143.680 ;
        RECT 110.360 139.600 110.620 139.920 ;
        RECT 110.420 134.480 110.560 139.600 ;
        RECT 110.360 134.160 110.620 134.480 ;
        RECT 110.880 134.140 111.020 154.560 ;
        RECT 111.340 134.140 111.480 170.880 ;
        RECT 112.660 169.180 112.920 169.500 ;
        RECT 111.740 168.840 112.000 169.160 ;
        RECT 111.800 166.440 111.940 168.840 ;
        RECT 112.200 166.460 112.460 166.780 ;
        RECT 111.740 166.120 112.000 166.440 ;
        RECT 112.260 166.100 112.400 166.460 ;
        RECT 112.200 165.780 112.460 166.100 ;
        RECT 111.740 163.060 112.000 163.380 ;
        RECT 111.800 158.700 111.940 163.060 ;
        RECT 112.260 159.300 112.400 165.780 ;
        RECT 112.720 163.720 112.860 169.180 ;
        RECT 113.120 168.160 113.380 168.480 ;
        RECT 113.180 164.740 113.320 168.160 ;
        RECT 113.120 164.420 113.380 164.740 ;
        RECT 113.180 163.720 113.320 164.420 ;
        RECT 112.660 163.400 112.920 163.720 ;
        RECT 113.120 163.400 113.380 163.720 ;
        RECT 112.720 161.000 112.860 163.400 ;
        RECT 112.660 160.680 112.920 161.000 ;
        RECT 112.200 158.980 112.460 159.300 ;
        RECT 111.800 158.560 112.400 158.700 ;
        RECT 111.740 157.960 112.000 158.280 ;
        RECT 111.800 156.580 111.940 157.960 ;
        RECT 112.260 157.940 112.400 158.560 ;
        RECT 112.200 157.620 112.460 157.940 ;
        RECT 111.740 156.260 112.000 156.580 ;
        RECT 112.260 152.160 112.400 157.620 ;
        RECT 113.180 155.900 113.320 163.400 ;
        RECT 113.640 163.380 113.780 170.880 ;
        RECT 114.560 169.160 114.700 171.220 ;
        RECT 117.260 170.880 117.520 171.200 ;
        RECT 117.320 169.500 117.460 170.880 ;
        RECT 117.260 169.180 117.520 169.500 ;
        RECT 114.500 168.840 114.760 169.160 ;
        RECT 114.040 165.440 114.300 165.760 ;
        RECT 113.580 163.060 113.840 163.380 ;
        RECT 114.100 161.340 114.240 165.440 ;
        RECT 114.040 161.020 114.300 161.340 ;
        RECT 113.120 155.580 113.380 155.900 ;
        RECT 114.560 153.520 114.700 168.840 ;
        RECT 117.320 162.020 117.460 169.180 ;
        RECT 116.340 161.700 116.600 162.020 ;
        RECT 117.260 161.700 117.520 162.020 ;
        RECT 114.500 153.200 114.760 153.520 ;
        RECT 116.400 153.180 116.540 161.700 ;
        RECT 119.160 161.340 119.300 172.580 ;
        RECT 121.400 171.560 121.660 171.880 ;
        RECT 124.620 171.560 124.880 171.880 ;
        RECT 121.460 170.180 121.600 171.560 ;
        RECT 121.800 170.345 123.680 170.715 ;
        RECT 121.400 169.860 121.660 170.180 ;
        RECT 119.560 166.800 119.820 167.120 ;
        RECT 119.620 162.020 119.760 166.800 ;
        RECT 124.680 166.780 124.820 171.560 ;
        RECT 127.830 171.365 128.110 171.735 ;
        RECT 127.900 169.160 128.040 171.365 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 127.840 168.840 128.100 169.160 ;
        RECT 124.620 166.460 124.880 166.780 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 121.400 165.440 121.660 165.760 ;
        RECT 121.460 162.020 121.600 165.440 ;
        RECT 121.800 164.905 123.680 165.275 ;
        RECT 124.680 164.060 124.820 166.460 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 124.620 163.740 124.880 164.060 ;
        RECT 123.700 163.400 123.960 163.720 ;
        RECT 119.560 161.700 119.820 162.020 ;
        RECT 121.400 161.700 121.660 162.020 ;
        RECT 123.760 161.680 123.900 163.400 ;
        RECT 123.700 161.360 123.960 161.680 ;
        RECT 119.100 161.020 119.360 161.340 ;
        RECT 120.940 161.020 121.200 161.340 ;
        RECT 116.800 160.000 117.060 160.320 ;
        RECT 116.860 158.620 117.000 160.000 ;
        RECT 121.000 159.300 121.140 161.020 ;
        RECT 121.800 159.465 123.680 159.835 ;
        RECT 120.940 158.980 121.200 159.300 ;
        RECT 116.800 158.300 117.060 158.620 ;
        RECT 117.720 155.240 117.980 155.560 ;
        RECT 116.340 152.860 116.600 153.180 ;
        RECT 115.880 152.180 116.140 152.500 ;
        RECT 112.200 151.840 112.460 152.160 ;
        RECT 111.740 149.460 112.000 149.780 ;
        RECT 111.800 145.020 111.940 149.460 ;
        RECT 114.040 149.120 114.300 149.440 ;
        RECT 113.120 147.420 113.380 147.740 ;
        RECT 112.200 147.080 112.460 147.400 ;
        RECT 111.740 144.700 112.000 145.020 ;
        RECT 112.260 144.930 112.400 147.080 ;
        RECT 112.660 144.930 112.920 145.020 ;
        RECT 112.260 144.790 112.920 144.930 ;
        RECT 112.660 144.700 112.920 144.790 ;
        RECT 111.800 143.740 111.940 144.700 ;
        RECT 113.180 144.590 113.320 147.420 ;
        RECT 114.100 146.720 114.240 149.120 ;
        RECT 115.940 148.420 116.080 152.180 ;
        RECT 116.800 150.710 117.060 150.800 ;
        RECT 117.780 150.710 117.920 155.240 ;
        RECT 121.800 154.025 123.680 154.395 ;
        RECT 119.560 152.520 119.820 152.840 ;
        RECT 118.180 151.840 118.440 152.160 ;
        RECT 118.240 150.800 118.380 151.840 ;
        RECT 116.800 150.570 117.920 150.710 ;
        RECT 116.800 150.480 117.060 150.570 ;
        RECT 115.880 148.100 116.140 148.420 ;
        RECT 117.780 147.650 117.920 150.570 ;
        RECT 118.180 150.480 118.440 150.800 ;
        RECT 117.780 147.510 118.380 147.650 ;
        RECT 117.720 146.740 117.980 147.060 ;
        RECT 114.040 146.400 114.300 146.720 ;
        RECT 117.260 146.400 117.520 146.720 ;
        RECT 117.320 145.700 117.460 146.400 ;
        RECT 117.260 145.380 117.520 145.700 ;
        RECT 117.780 144.680 117.920 146.740 ;
        RECT 113.580 144.590 113.840 144.680 ;
        RECT 113.180 144.450 113.840 144.590 ;
        RECT 111.800 143.600 112.860 143.740 ;
        RECT 111.740 142.660 112.000 142.980 ;
        RECT 110.820 133.820 111.080 134.140 ;
        RECT 111.280 133.820 111.540 134.140 ;
        RECT 110.360 132.800 110.620 133.120 ;
        RECT 111.280 132.800 111.540 133.120 ;
        RECT 109.900 131.780 110.160 132.100 ;
        RECT 106.800 129.545 108.680 129.915 ;
        RECT 104.840 129.060 105.100 129.380 ;
        RECT 106.220 129.060 106.480 129.380 ;
        RECT 106.220 128.380 106.480 128.700 ;
        RECT 105.300 128.040 105.560 128.360 ;
        RECT 105.360 125.640 105.500 128.040 ;
        RECT 105.300 125.320 105.560 125.640 ;
        RECT 105.300 122.600 105.560 122.920 ;
        RECT 105.360 120.540 105.500 122.600 ;
        RECT 105.300 120.220 105.560 120.540 ;
        RECT 106.280 119.860 106.420 128.380 ;
        RECT 109.440 128.040 109.700 128.360 ;
        RECT 106.800 124.105 108.680 124.475 ;
        RECT 109.500 120.540 109.640 128.040 ;
        RECT 109.440 120.220 109.700 120.540 ;
        RECT 106.220 119.540 106.480 119.860 ;
        RECT 105.760 119.200 106.020 119.520 ;
        RECT 108.980 119.200 109.240 119.520 ;
        RECT 105.820 118.160 105.960 119.200 ;
        RECT 106.800 118.665 108.680 119.035 ;
        RECT 105.760 117.840 106.020 118.160 ;
        RECT 109.040 114.760 109.180 119.200 ;
        RECT 109.500 114.760 109.640 120.220 ;
        RECT 109.900 117.500 110.160 117.820 ;
        RECT 109.960 115.780 110.100 117.500 ;
        RECT 109.900 115.460 110.160 115.780 ;
        RECT 108.980 114.440 109.240 114.760 ;
        RECT 109.440 114.440 109.700 114.760 ;
        RECT 106.800 113.225 108.680 113.595 ;
        RECT 104.380 111.720 104.640 112.040 ;
        RECT 110.420 109.320 110.560 132.800 ;
        RECT 110.820 130.760 111.080 131.080 ;
        RECT 110.880 128.700 111.020 130.760 ;
        RECT 111.340 129.380 111.480 132.800 ;
        RECT 111.280 129.060 111.540 129.380 ;
        RECT 111.800 128.780 111.940 142.660 ;
        RECT 112.200 139.600 112.460 139.920 ;
        RECT 112.260 134.480 112.400 139.600 ;
        RECT 112.720 139.580 112.860 143.600 ;
        RECT 113.180 142.300 113.320 144.450 ;
        RECT 113.580 144.360 113.840 144.450 ;
        RECT 117.720 144.360 117.980 144.680 ;
        RECT 113.120 141.980 113.380 142.300 ;
        RECT 112.660 139.260 112.920 139.580 ;
        RECT 112.660 138.580 112.920 138.900 ;
        RECT 112.720 136.520 112.860 138.580 ;
        RECT 113.180 137.200 113.320 141.980 ;
        RECT 117.780 141.960 117.920 144.360 ;
        RECT 117.720 141.640 117.980 141.960 ;
        RECT 117.260 140.960 117.520 141.280 ;
        RECT 117.320 139.920 117.460 140.960 ;
        RECT 117.260 139.600 117.520 139.920 ;
        RECT 115.880 139.260 116.140 139.580 ;
        RECT 113.120 136.880 113.380 137.200 ;
        RECT 112.660 136.200 112.920 136.520 ;
        RECT 115.940 136.180 116.080 139.260 ;
        RECT 115.880 135.860 116.140 136.180 ;
        RECT 113.120 135.520 113.380 135.840 ;
        RECT 112.200 134.160 112.460 134.480 ;
        RECT 113.180 134.140 113.320 135.520 ;
        RECT 113.120 133.820 113.380 134.140 ;
        RECT 118.240 131.760 118.380 147.510 ;
        RECT 119.620 145.020 119.760 152.520 ;
        RECT 123.240 151.840 123.500 152.160 ;
        RECT 123.300 150.800 123.440 151.840 ;
        RECT 123.240 150.480 123.500 150.800 ;
        RECT 126.000 149.800 126.260 150.120 ;
        RECT 121.800 148.585 123.680 148.955 ;
        RECT 126.060 147.400 126.200 149.800 ;
        RECT 123.700 147.080 123.960 147.400 ;
        RECT 126.000 147.080 126.260 147.400 ;
        RECT 120.020 146.740 120.280 147.060 ;
        RECT 120.080 145.700 120.220 146.740 ;
        RECT 123.760 145.700 123.900 147.080 ;
        RECT 120.020 145.380 120.280 145.700 ;
        RECT 123.700 145.380 123.960 145.700 ;
        RECT 119.560 144.700 119.820 145.020 ;
        RECT 119.620 141.960 119.760 144.700 ;
        RECT 121.800 143.145 123.680 143.515 ;
        RECT 119.560 141.700 119.820 141.960 ;
        RECT 119.560 141.640 120.220 141.700 ;
        RECT 119.620 141.560 120.220 141.640 ;
        RECT 119.560 140.960 119.820 141.280 ;
        RECT 119.620 137.540 119.760 140.960 ;
        RECT 120.080 138.900 120.220 141.560 ;
        RECT 120.480 140.960 120.740 141.280 ;
        RECT 120.540 139.920 120.680 140.960 ;
        RECT 120.480 139.600 120.740 139.920 ;
        RECT 124.160 139.260 124.420 139.580 ;
        RECT 120.020 138.580 120.280 138.900 ;
        RECT 121.400 138.240 121.660 138.560 ;
        RECT 119.560 137.220 119.820 137.540 ;
        RECT 121.460 136.860 121.600 138.240 ;
        RECT 121.800 137.705 123.680 138.075 ;
        RECT 124.220 137.540 124.360 139.260 ;
        RECT 126.060 139.240 126.200 147.080 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 126.000 138.920 126.260 139.240 ;
        RECT 124.620 138.240 124.880 138.560 ;
        RECT 124.160 137.220 124.420 137.540 ;
        RECT 121.400 136.540 121.660 136.860 ;
        RECT 120.940 136.200 121.200 136.520 ;
        RECT 121.000 134.820 121.140 136.200 ;
        RECT 120.940 134.500 121.200 134.820 ;
        RECT 121.800 132.265 123.680 132.635 ;
        RECT 118.180 131.440 118.440 131.760 ;
        RECT 112.200 130.760 112.460 131.080 ;
        RECT 110.820 128.380 111.080 128.700 ;
        RECT 111.340 128.640 111.940 128.780 ;
        RECT 110.820 109.680 111.080 110.000 ;
        RECT 94.720 109.000 94.980 109.320 ;
        RECT 99.780 109.000 100.040 109.320 ;
        RECT 103.460 109.000 103.720 109.320 ;
        RECT 110.360 109.000 110.620 109.320 ;
        RECT 102.540 108.660 102.800 108.980 ;
        RECT 87.820 108.320 88.080 108.640 ;
        RECT 92.880 108.320 93.140 108.640 ;
        RECT 97.940 108.320 98.200 108.640 ;
        RECT 99.780 108.320 100.040 108.640 ;
        RECT 86.900 106.620 87.160 106.940 ;
        RECT 80.000 106.280 80.260 106.600 ;
        RECT 86.440 106.280 86.700 106.600 ;
        RECT 79.540 103.560 79.800 103.880 ;
        RECT 74.020 103.220 74.280 103.540 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 56.070 89.190 56.350 89.210 ;
        RECT 55.530 88.660 56.750 89.190 ;
        RECT 62.050 88.870 62.330 89.210 ;
        RECT 37.680 86.810 39.070 88.520 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 54.760 88.520 56.750 88.660 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 88.520 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 74.080 89.210 74.220 103.220 ;
        RECT 76.800 102.345 78.680 102.715 ;
        RECT 80.060 89.210 80.200 106.280 ;
        RECT 86.500 104.220 86.640 106.280 ;
        RECT 86.440 103.900 86.700 104.220 ;
        RECT 87.880 103.540 88.020 108.320 ;
        RECT 92.940 107.280 93.080 108.320 ;
        RECT 93.800 107.300 94.060 107.620 ;
        RECT 92.880 106.960 93.140 107.280 ;
        RECT 88.280 105.600 88.540 105.920 ;
        RECT 88.340 104.220 88.480 105.600 ;
        RECT 91.800 105.065 93.680 105.435 ;
        RECT 88.280 103.900 88.540 104.220 ;
        RECT 86.900 103.220 87.160 103.540 ;
        RECT 87.820 103.220 88.080 103.540 ;
        RECT 74.010 88.160 74.290 89.210 ;
        RECT 79.990 88.180 80.270 89.210 ;
        RECT 85.970 88.660 86.250 89.210 ;
        RECT 86.960 88.660 87.100 103.220 ;
        RECT 91.800 99.625 93.680 99.995 ;
        RECT 85.970 88.520 87.100 88.660 ;
        RECT 91.950 88.660 92.230 89.210 ;
        RECT 93.860 88.660 94.000 107.300 ;
        RECT 98.000 107.280 98.140 108.320 ;
        RECT 97.940 106.960 98.200 107.280 ;
        RECT 99.320 106.280 99.580 106.600 ;
        RECT 97.480 105.600 97.740 105.920 ;
        RECT 97.540 101.840 97.680 105.600 ;
        RECT 99.380 104.220 99.520 106.280 ;
        RECT 99.320 103.900 99.580 104.220 ;
        RECT 97.480 101.520 97.740 101.840 ;
        RECT 99.380 101.160 99.520 103.900 ;
        RECT 99.840 101.840 99.980 108.320 ;
        RECT 102.600 106.940 102.740 108.660 ;
        RECT 109.440 108.320 109.700 108.640 ;
        RECT 106.800 107.785 108.680 108.155 ;
        RECT 108.980 107.300 109.240 107.620 ;
        RECT 102.540 106.620 102.800 106.940 ;
        RECT 104.380 105.600 104.640 105.920 ;
        RECT 104.440 103.540 104.580 105.600 ;
        RECT 103.920 103.220 104.180 103.540 ;
        RECT 104.380 103.220 104.640 103.540 ;
        RECT 99.780 101.520 100.040 101.840 ;
        RECT 97.940 100.840 98.200 101.160 ;
        RECT 99.320 100.840 99.580 101.160 ;
        RECT 98.000 89.210 98.140 100.840 ;
        RECT 103.980 89.210 104.120 103.220 ;
        RECT 106.800 102.345 108.680 102.715 ;
        RECT 109.040 98.180 109.180 107.300 ;
        RECT 109.500 107.280 109.640 108.320 ;
        RECT 109.440 106.960 109.700 107.280 ;
        RECT 110.880 104.220 111.020 109.680 ;
        RECT 111.340 109.320 111.480 128.640 ;
        RECT 112.260 125.550 112.400 130.760 ;
        RECT 118.240 128.700 118.380 131.440 ;
        RECT 113.120 128.380 113.380 128.700 ;
        RECT 118.180 128.380 118.440 128.700 ;
        RECT 112.260 125.410 112.860 125.550 ;
        RECT 112.720 123.260 112.860 125.410 ;
        RECT 113.180 124.960 113.320 128.380 ;
        RECT 114.960 128.040 115.220 128.360 ;
        RECT 115.020 126.660 115.160 128.040 ;
        RECT 114.960 126.340 115.220 126.660 ;
        RECT 113.580 125.660 113.840 125.980 ;
        RECT 113.120 124.640 113.380 124.960 ;
        RECT 113.180 123.600 113.320 124.640 ;
        RECT 113.120 123.280 113.380 123.600 ;
        RECT 112.660 122.940 112.920 123.260 ;
        RECT 111.740 119.200 112.000 119.520 ;
        RECT 111.800 117.820 111.940 119.200 ;
        RECT 111.740 117.500 112.000 117.820 ;
        RECT 111.800 113.060 111.940 117.500 ;
        RECT 112.720 115.100 112.860 122.940 ;
        RECT 113.640 122.920 113.780 125.660 ;
        RECT 113.580 122.830 113.840 122.920 ;
        RECT 113.180 122.690 113.840 122.830 ;
        RECT 113.180 115.440 113.320 122.690 ;
        RECT 113.580 122.600 113.840 122.690 ;
        RECT 116.340 119.880 116.600 120.200 ;
        RECT 118.240 120.110 118.380 128.380 ;
        RECT 118.640 127.360 118.900 127.680 ;
        RECT 120.480 127.360 120.740 127.680 ;
        RECT 118.700 125.300 118.840 127.360 ;
        RECT 120.540 125.980 120.680 127.360 ;
        RECT 121.800 126.825 123.680 127.195 ;
        RECT 120.480 125.660 120.740 125.980 ;
        RECT 124.680 125.640 124.820 138.240 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 124.620 125.320 124.880 125.640 ;
        RECT 118.640 124.980 118.900 125.300 ;
        RECT 119.100 123.280 119.360 123.600 ;
        RECT 119.160 121.220 119.300 123.280 ;
        RECT 124.680 123.260 124.820 125.320 ;
        RECT 124.620 122.940 124.880 123.260 ;
        RECT 121.400 122.600 121.660 122.920 ;
        RECT 120.480 121.920 120.740 122.240 ;
        RECT 119.100 120.900 119.360 121.220 ;
        RECT 120.540 120.200 120.680 121.920 ;
        RECT 121.460 121.220 121.600 122.600 ;
        RECT 121.800 121.385 123.680 121.755 ;
        RECT 121.400 120.900 121.660 121.220 ;
        RECT 118.640 120.110 118.900 120.200 ;
        RECT 118.240 119.970 118.900 120.110 ;
        RECT 113.580 119.540 113.840 119.860 ;
        RECT 113.640 118.500 113.780 119.540 ;
        RECT 116.400 118.500 116.540 119.880 ;
        RECT 113.580 118.180 113.840 118.500 ;
        RECT 116.340 118.180 116.600 118.500 ;
        RECT 118.240 118.160 118.380 119.970 ;
        RECT 118.640 119.880 118.900 119.970 ;
        RECT 120.480 119.880 120.740 120.200 ;
        RECT 118.180 117.840 118.440 118.160 ;
        RECT 115.420 117.500 115.680 117.820 ;
        RECT 115.480 115.780 115.620 117.500 ;
        RECT 121.800 115.945 123.680 116.315 ;
        RECT 115.420 115.460 115.680 115.780 ;
        RECT 113.120 115.120 113.380 115.440 ;
        RECT 112.660 114.780 112.920 115.100 ;
        RECT 121.860 113.760 122.120 114.080 ;
        RECT 111.740 112.740 112.000 113.060 ;
        RECT 117.260 112.740 117.520 113.060 ;
        RECT 111.800 110.000 111.940 112.740 ;
        RECT 111.740 109.680 112.000 110.000 ;
        RECT 111.280 109.000 111.540 109.320 ;
        RECT 111.280 108.320 111.540 108.640 ;
        RECT 111.340 107.280 111.480 108.320 ;
        RECT 111.280 106.960 111.540 107.280 ;
        RECT 111.800 107.020 111.940 109.680 ;
        RECT 114.040 108.320 114.300 108.640 ;
        RECT 116.340 108.320 116.600 108.640 ;
        RECT 111.800 106.880 112.400 107.020 ;
        RECT 112.260 106.600 112.400 106.880 ;
        RECT 112.200 106.280 112.460 106.600 ;
        RECT 112.260 104.220 112.400 106.280 ;
        RECT 114.100 104.220 114.240 108.320 ;
        RECT 110.820 103.900 111.080 104.220 ;
        RECT 112.200 103.900 112.460 104.220 ;
        RECT 114.040 103.900 114.300 104.220 ;
        RECT 115.880 103.900 116.140 104.220 ;
        RECT 109.040 98.040 110.100 98.180 ;
        RECT 109.960 89.290 110.100 98.040 ;
        RECT 115.940 89.570 116.080 103.900 ;
        RECT 116.400 103.540 116.540 108.320 ;
        RECT 117.320 107.280 117.460 112.740 ;
        RECT 119.100 112.400 119.360 112.720 ;
        RECT 119.160 109.660 119.300 112.400 ;
        RECT 121.920 112.380 122.060 113.760 ;
        RECT 119.560 112.060 119.820 112.380 ;
        RECT 121.860 112.060 122.120 112.380 ;
        RECT 119.100 109.340 119.360 109.660 ;
        RECT 119.100 108.550 119.360 108.640 ;
        RECT 119.620 108.550 119.760 112.060 ;
        RECT 120.020 111.720 120.280 112.040 ;
        RECT 120.080 108.980 120.220 111.720 ;
        RECT 121.800 110.505 123.680 110.875 ;
        RECT 120.020 108.660 120.280 108.980 ;
        RECT 127.840 108.660 128.100 108.980 ;
        RECT 119.100 108.410 119.760 108.550 ;
        RECT 119.100 108.320 119.360 108.410 ;
        RECT 117.260 106.960 117.520 107.280 ;
        RECT 116.340 103.220 116.600 103.540 ;
        RECT 119.620 101.500 119.760 108.410 ;
        RECT 120.020 106.960 120.280 107.280 ;
        RECT 120.080 102.180 120.220 106.960 ;
        RECT 120.940 106.280 121.200 106.600 ;
        RECT 120.020 101.860 120.280 102.180 ;
        RECT 119.560 101.180 119.820 101.500 ;
        RECT 121.000 98.860 121.140 106.280 ;
        RECT 125.990 106.085 126.270 106.455 ;
        RECT 121.800 105.065 123.680 105.435 ;
        RECT 126.060 103.880 126.200 106.085 ;
        RECT 126.000 103.560 126.260 103.880 ;
        RECT 121.800 99.625 123.680 99.995 ;
        RECT 121.000 98.720 122.060 98.860 ;
        RECT 121.920 89.570 122.060 98.720 ;
        RECT 91.950 88.520 94.000 88.660 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 85.970 87.970 86.250 88.520 ;
        RECT 91.950 88.320 92.230 88.520 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.930 88.240 98.210 89.210 ;
        RECT 103.910 88.610 104.190 89.210 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 127.900 89.380 128.040 108.660 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 16.750 211.165 18.730 211.495 ;
        RECT 46.750 211.165 48.730 211.495 ;
        RECT 76.750 211.165 78.730 211.495 ;
        RECT 106.750 211.165 108.730 211.495 ;
        RECT 31.750 208.445 33.730 208.775 ;
        RECT 61.750 208.445 63.730 208.775 ;
        RECT 91.750 208.445 93.730 208.775 ;
        RECT 121.750 208.445 123.730 208.775 ;
        RECT 16.750 205.725 18.730 206.055 ;
        RECT 46.750 205.725 48.730 206.055 ;
        RECT 76.750 205.725 78.730 206.055 ;
        RECT 106.750 205.725 108.730 206.055 ;
        RECT 31.750 203.005 33.730 203.335 ;
        RECT 61.750 203.005 63.730 203.335 ;
        RECT 91.750 203.005 93.730 203.335 ;
        RECT 121.750 203.005 123.730 203.335 ;
        RECT 16.750 200.285 18.730 200.615 ;
        RECT 46.750 200.285 48.730 200.615 ;
        RECT 76.750 200.285 78.730 200.615 ;
        RECT 106.750 200.285 108.730 200.615 ;
        RECT 31.750 197.565 33.730 197.895 ;
        RECT 61.750 197.565 63.730 197.895 ;
        RECT 91.750 197.565 93.730 197.895 ;
        RECT 121.750 197.565 123.730 197.895 ;
        RECT 16.750 194.845 18.730 195.175 ;
        RECT 46.750 194.845 48.730 195.175 ;
        RECT 76.750 194.845 78.730 195.175 ;
        RECT 106.750 194.845 108.730 195.175 ;
        RECT 31.750 192.125 33.730 192.455 ;
        RECT 61.750 192.125 63.730 192.455 ;
        RECT 91.750 192.125 93.730 192.455 ;
        RECT 121.750 192.125 123.730 192.455 ;
        RECT 16.750 189.405 18.730 189.735 ;
        RECT 46.750 189.405 48.730 189.735 ;
        RECT 76.750 189.405 78.730 189.735 ;
        RECT 106.750 189.405 108.730 189.735 ;
        RECT 44.290 188.020 44.670 188.030 ;
        RECT 55.585 188.020 55.915 188.035 ;
        RECT 44.290 187.720 55.915 188.020 ;
        RECT 44.290 187.710 44.670 187.720 ;
        RECT 55.585 187.705 55.915 187.720 ;
        RECT 94.685 188.020 95.015 188.035 ;
        RECT 98.570 188.020 98.950 188.030 ;
        RECT 94.685 187.720 98.950 188.020 ;
        RECT 94.685 187.705 95.015 187.720 ;
        RECT 98.570 187.710 98.950 187.720 ;
        RECT 31.750 186.685 33.730 187.015 ;
        RECT 61.750 186.685 63.730 187.015 ;
        RECT 91.750 186.685 93.730 187.015 ;
        RECT 121.750 186.685 123.730 187.015 ;
        RECT 16.750 183.965 18.730 184.295 ;
        RECT 46.750 183.965 48.730 184.295 ;
        RECT 76.750 183.965 78.730 184.295 ;
        RECT 106.750 183.965 108.730 184.295 ;
        RECT 31.750 181.245 33.730 181.575 ;
        RECT 61.750 181.245 63.730 181.575 ;
        RECT 91.750 181.245 93.730 181.575 ;
        RECT 121.750 181.245 123.730 181.575 ;
        RECT 40.405 179.860 40.735 179.875 ;
        RECT 41.785 179.860 42.115 179.875 ;
        RECT 67.545 179.860 67.875 179.875 ;
        RECT 40.405 179.560 67.875 179.860 ;
        RECT 40.405 179.545 40.735 179.560 ;
        RECT 41.785 179.545 42.115 179.560 ;
        RECT 67.545 179.545 67.875 179.560 ;
        RECT 78.585 179.860 78.915 179.875 ;
        RECT 85.025 179.860 85.355 179.875 ;
        RECT 78.585 179.560 85.355 179.860 ;
        RECT 78.585 179.545 78.915 179.560 ;
        RECT 85.025 179.545 85.355 179.560 ;
        RECT 16.750 178.525 18.730 178.855 ;
        RECT 46.750 178.525 48.730 178.855 ;
        RECT 76.750 178.525 78.730 178.855 ;
        RECT 106.750 178.525 108.730 178.855 ;
        RECT 66.165 177.820 66.495 177.835 ;
        RECT 70.305 177.820 70.635 177.835 ;
        RECT 72.605 177.820 72.935 177.835 ;
        RECT 66.165 177.520 72.935 177.820 ;
        RECT 66.165 177.505 66.495 177.520 ;
        RECT 70.305 177.505 70.635 177.520 ;
        RECT 72.605 177.505 72.935 177.520 ;
        RECT 71.685 177.140 72.015 177.155 ;
        RECT 78.125 177.140 78.455 177.155 ;
        RECT 71.685 176.840 78.455 177.140 ;
        RECT 71.685 176.825 72.015 176.840 ;
        RECT 78.125 176.825 78.455 176.840 ;
        RECT 31.750 175.805 33.730 176.135 ;
        RECT 61.750 175.805 63.730 176.135 ;
        RECT 91.750 175.805 93.730 176.135 ;
        RECT 121.750 175.805 123.730 176.135 ;
        RECT 39.945 175.100 40.275 175.115 ;
        RECT 65.245 175.100 65.575 175.115 ;
        RECT 39.945 174.800 65.575 175.100 ;
        RECT 39.945 174.785 40.275 174.800 ;
        RECT 65.245 174.785 65.575 174.800 ;
        RECT 54.665 174.420 54.995 174.435 ;
        RECT 62.945 174.420 63.275 174.435 ;
        RECT 54.665 174.120 63.275 174.420 ;
        RECT 54.665 174.105 54.995 174.120 ;
        RECT 62.945 174.105 63.275 174.120 ;
        RECT 16.750 173.085 18.730 173.415 ;
        RECT 46.750 173.085 48.730 173.415 ;
        RECT 76.750 173.085 78.730 173.415 ;
        RECT 106.750 173.085 108.730 173.415 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 127.805 171.700 128.135 171.715 ;
        RECT 129.030 171.700 134.930 172.500 ;
        RECT 127.805 171.400 134.930 171.700 ;
        RECT 127.805 171.385 128.135 171.400 ;
        RECT 31.750 170.365 33.730 170.695 ;
        RECT 61.750 170.365 63.730 170.695 ;
        RECT 91.750 170.365 93.730 170.695 ;
        RECT 121.750 170.365 123.730 170.695 ;
        RECT 129.030 170.130 134.930 171.400 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 44.085 169.670 44.415 169.675 ;
        RECT 44.085 169.660 44.670 169.670 ;
        RECT 43.860 169.360 44.670 169.660 ;
        RECT 44.085 169.350 44.670 169.360 ;
        RECT 44.085 169.345 44.415 169.350 ;
        RECT 16.750 167.645 18.730 167.975 ;
        RECT 46.750 167.645 48.730 167.975 ;
        RECT 76.750 167.645 78.730 167.975 ;
        RECT 106.750 167.645 108.730 167.975 ;
        RECT 31.750 164.925 33.730 165.255 ;
        RECT 61.750 164.925 63.730 165.255 ;
        RECT 91.750 164.925 93.730 165.255 ;
        RECT 121.750 164.925 123.730 165.255 ;
        RECT 94.890 164.220 95.270 164.230 ;
        RECT 98.570 164.220 98.950 164.230 ;
        RECT 101.125 164.220 101.455 164.235 ;
        RECT 94.890 163.920 101.455 164.220 ;
        RECT 94.890 163.910 95.270 163.920 ;
        RECT 98.570 163.910 98.950 163.920 ;
        RECT 101.125 163.905 101.455 163.920 ;
        RECT 16.750 162.205 18.730 162.535 ;
        RECT 46.750 162.205 48.730 162.535 ;
        RECT 76.750 162.205 78.730 162.535 ;
        RECT 106.750 162.205 108.730 162.535 ;
        RECT 31.750 159.485 33.730 159.815 ;
        RECT 61.750 159.485 63.730 159.815 ;
        RECT 91.750 159.485 93.730 159.815 ;
        RECT 121.750 159.485 123.730 159.815 ;
        RECT 79.965 159.460 80.295 159.475 ;
        RECT 81.345 159.460 81.675 159.475 ;
        RECT 79.965 159.160 81.675 159.460 ;
        RECT 79.965 159.145 80.295 159.160 ;
        RECT 81.345 159.145 81.675 159.160 ;
        RECT 68.005 158.780 68.335 158.795 ;
        RECT 71.685 158.780 72.015 158.795 ;
        RECT 84.565 158.780 84.895 158.795 ;
        RECT 68.005 158.480 84.895 158.780 ;
        RECT 68.005 158.465 68.335 158.480 ;
        RECT 71.685 158.465 72.015 158.480 ;
        RECT 84.565 158.465 84.895 158.480 ;
        RECT 16.750 156.765 18.730 157.095 ;
        RECT 46.750 156.765 48.730 157.095 ;
        RECT 76.750 156.765 78.730 157.095 ;
        RECT 106.750 156.765 108.730 157.095 ;
        RECT 73.065 156.740 73.395 156.755 ;
        RECT 75.365 156.740 75.695 156.755 ;
        RECT 73.065 156.440 75.695 156.740 ;
        RECT 73.065 156.425 73.395 156.440 ;
        RECT 75.365 156.425 75.695 156.440 ;
        RECT 41.785 156.060 42.115 156.075 ;
        RECT 43.165 156.060 43.495 156.075 ;
        RECT 94.890 156.060 95.270 156.070 ;
        RECT 41.785 155.760 43.495 156.060 ;
        RECT 41.785 155.745 42.115 155.760 ;
        RECT 43.165 155.745 43.495 155.760 ;
        RECT 71.010 155.760 95.270 156.060 ;
        RECT 44.290 155.380 44.670 155.390 ;
        RECT 65.705 155.380 66.035 155.395 ;
        RECT 71.010 155.380 71.310 155.760 ;
        RECT 94.890 155.750 95.270 155.760 ;
        RECT 44.290 155.080 71.310 155.380 ;
        RECT 74.445 155.380 74.775 155.395 ;
        RECT 112.370 155.380 112.750 155.390 ;
        RECT 74.445 155.080 112.750 155.380 ;
        RECT 44.290 155.070 44.670 155.080 ;
        RECT 65.705 155.065 66.035 155.080 ;
        RECT 74.445 155.065 74.775 155.080 ;
        RECT 112.370 155.070 112.750 155.080 ;
        RECT 31.750 154.045 33.730 154.375 ;
        RECT 61.750 154.045 63.730 154.375 ;
        RECT 91.750 154.045 93.730 154.375 ;
        RECT 121.750 154.045 123.730 154.375 ;
        RECT 44.545 152.660 44.875 152.675 ;
        RECT 68.005 152.660 68.335 152.675 ;
        RECT 44.545 152.360 68.335 152.660 ;
        RECT 44.545 152.345 44.875 152.360 ;
        RECT 68.005 152.345 68.335 152.360 ;
        RECT 16.750 151.325 18.730 151.655 ;
        RECT 46.750 151.325 48.730 151.655 ;
        RECT 76.750 151.325 78.730 151.655 ;
        RECT 106.750 151.325 108.730 151.655 ;
        RECT 87.785 150.620 88.115 150.635 ;
        RECT 99.285 150.620 99.615 150.635 ;
        RECT 107.565 150.620 107.895 150.635 ;
        RECT 87.785 150.320 107.895 150.620 ;
        RECT 87.785 150.305 88.115 150.320 ;
        RECT 99.285 150.305 99.615 150.320 ;
        RECT 107.565 150.305 107.895 150.320 ;
        RECT 31.750 148.605 33.730 148.935 ;
        RECT 61.750 148.605 63.730 148.935 ;
        RECT 91.750 148.605 93.730 148.935 ;
        RECT 121.750 148.605 123.730 148.935 ;
        RECT 16.750 145.885 18.730 146.215 ;
        RECT 46.750 145.885 48.730 146.215 ;
        RECT 76.750 145.885 78.730 146.215 ;
        RECT 106.750 145.885 108.730 146.215 ;
        RECT 31.750 143.165 33.730 143.495 ;
        RECT 61.750 143.165 63.730 143.495 ;
        RECT 91.750 143.165 93.730 143.495 ;
        RECT 121.750 143.165 123.730 143.495 ;
        RECT 16.750 140.445 18.730 140.775 ;
        RECT 46.750 140.445 48.730 140.775 ;
        RECT 76.750 140.445 78.730 140.775 ;
        RECT 106.750 140.445 108.730 140.775 ;
        RECT 132.510 139.210 135.210 140.035 ;
        RECT 112.370 139.060 112.750 139.070 ;
        RECT 131.260 139.060 135.210 139.210 ;
        RECT 112.370 138.760 135.210 139.060 ;
        RECT 112.370 138.750 112.750 138.760 ;
        RECT 131.260 138.610 135.210 138.760 ;
        RECT 132.510 138.165 135.210 138.610 ;
        RECT 31.750 137.725 33.730 138.055 ;
        RECT 61.750 137.725 63.730 138.055 ;
        RECT 91.750 137.725 93.730 138.055 ;
        RECT 121.750 137.725 123.730 138.055 ;
        RECT 16.750 135.005 18.730 135.335 ;
        RECT 46.750 135.005 48.730 135.335 ;
        RECT 76.750 135.005 78.730 135.335 ;
        RECT 106.750 135.005 108.730 135.335 ;
        RECT 99.285 134.300 99.615 134.315 ;
        RECT 108.025 134.300 108.355 134.315 ;
        RECT 99.285 134.000 108.355 134.300 ;
        RECT 99.285 133.985 99.615 134.000 ;
        RECT 108.025 133.985 108.355 134.000 ;
        RECT 31.750 132.285 33.730 132.615 ;
        RECT 61.750 132.285 63.730 132.615 ;
        RECT 91.750 132.285 93.730 132.615 ;
        RECT 121.750 132.285 123.730 132.615 ;
        RECT 44.290 132.260 44.670 132.270 ;
        RECT 49.145 132.260 49.475 132.275 ;
        RECT 44.290 131.960 49.475 132.260 ;
        RECT 44.290 131.950 44.670 131.960 ;
        RECT 49.145 131.945 49.475 131.960 ;
        RECT 16.750 129.565 18.730 129.895 ;
        RECT 46.750 129.565 48.730 129.895 ;
        RECT 76.750 129.565 78.730 129.895 ;
        RECT 106.750 129.565 108.730 129.895 ;
        RECT 94.890 129.540 95.270 129.550 ;
        RECT 95.605 129.540 95.935 129.555 ;
        RECT 94.890 129.240 95.935 129.540 ;
        RECT 94.890 129.230 95.270 129.240 ;
        RECT 95.605 129.225 95.935 129.240 ;
        RECT 31.750 126.845 33.730 127.175 ;
        RECT 61.750 126.845 63.730 127.175 ;
        RECT 91.750 126.845 93.730 127.175 ;
        RECT 121.750 126.845 123.730 127.175 ;
        RECT 16.750 124.125 18.730 124.455 ;
        RECT 46.750 124.125 48.730 124.455 ;
        RECT 76.750 124.125 78.730 124.455 ;
        RECT 106.750 124.125 108.730 124.455 ;
        RECT 31.750 121.405 33.730 121.735 ;
        RECT 61.750 121.405 63.730 121.735 ;
        RECT 91.750 121.405 93.730 121.735 ;
        RECT 121.750 121.405 123.730 121.735 ;
        RECT 16.750 118.685 18.730 119.015 ;
        RECT 46.750 118.685 48.730 119.015 ;
        RECT 76.750 118.685 78.730 119.015 ;
        RECT 106.750 118.685 108.730 119.015 ;
        RECT 31.750 115.965 33.730 116.295 ;
        RECT 61.750 115.965 63.730 116.295 ;
        RECT 91.750 115.965 93.730 116.295 ;
        RECT 121.750 115.965 123.730 116.295 ;
        RECT 16.750 113.245 18.730 113.575 ;
        RECT 46.750 113.245 48.730 113.575 ;
        RECT 76.750 113.245 78.730 113.575 ;
        RECT 106.750 113.245 108.730 113.575 ;
        RECT 92.845 113.220 93.175 113.235 ;
        RECT 94.890 113.220 95.270 113.230 ;
        RECT 92.845 112.920 95.270 113.220 ;
        RECT 92.845 112.905 93.175 112.920 ;
        RECT 94.890 112.910 95.270 112.920 ;
        RECT 31.750 110.525 33.730 110.855 ;
        RECT 61.750 110.525 63.730 110.855 ;
        RECT 91.750 110.525 93.730 110.855 ;
        RECT 121.750 110.525 123.730 110.855 ;
        RECT 16.750 107.805 18.730 108.135 ;
        RECT 46.750 107.805 48.730 108.135 ;
        RECT 76.750 107.805 78.730 108.135 ;
        RECT 106.750 107.805 108.730 108.135 ;
        RECT 129.700 106.570 133.210 106.625 ;
        RECT 125.965 106.420 126.295 106.435 ;
        RECT 129.700 106.420 133.260 106.570 ;
        RECT 125.965 106.120 133.260 106.420 ;
        RECT 125.965 106.105 126.295 106.120 ;
        RECT 129.700 105.970 133.260 106.120 ;
        RECT 129.700 105.605 133.210 105.970 ;
        RECT 31.750 105.085 33.730 105.415 ;
        RECT 61.750 105.085 63.730 105.415 ;
        RECT 91.750 105.085 93.730 105.415 ;
        RECT 121.750 105.085 123.730 105.415 ;
        RECT 16.750 102.365 18.730 102.695 ;
        RECT 46.750 102.365 48.730 102.695 ;
        RECT 76.750 102.365 78.730 102.695 ;
        RECT 106.750 102.365 108.730 102.695 ;
        RECT 31.750 99.645 33.730 99.975 ;
        RECT 61.750 99.645 63.730 99.975 ;
        RECT 91.750 99.645 93.730 99.975 ;
        RECT 121.750 99.645 123.730 99.975 ;
        RECT 1.040 98.100 11.400 98.110 ;
        RECT 1.040 97.980 11.420 98.100 ;
        RECT 0.970 96.160 11.420 97.980 ;
        RECT 0.970 96.140 3.030 96.160 ;
        RECT 9.420 96.100 11.420 96.160 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.740 99.570 18.740 211.570 ;
        RECT 31.740 101.605 33.740 211.570 ;
        RECT 44.315 187.705 44.645 188.035 ;
        RECT 44.330 169.675 44.630 187.705 ;
        RECT 44.315 169.345 44.645 169.675 ;
        RECT 44.330 155.395 44.630 169.345 ;
        RECT 44.315 155.065 44.645 155.395 ;
        RECT 44.330 132.275 44.630 155.065 ;
        RECT 44.315 131.945 44.645 132.275 ;
        RECT 31.740 99.570 33.770 101.605 ;
        RECT 46.740 99.570 48.740 211.570 ;
        RECT 61.740 99.570 63.740 211.570 ;
        RECT 76.740 99.570 78.740 211.570 ;
        RECT 91.740 99.570 93.740 211.570 ;
        RECT 98.595 187.705 98.925 188.035 ;
        RECT 98.610 164.235 98.910 187.705 ;
        RECT 94.915 163.905 95.245 164.235 ;
        RECT 98.595 163.905 98.925 164.235 ;
        RECT 94.930 156.075 95.230 163.905 ;
        RECT 94.915 155.745 95.245 156.075 ;
        RECT 94.930 129.555 95.230 155.745 ;
        RECT 94.915 129.225 95.245 129.555 ;
        RECT 94.930 113.235 95.230 129.225 ;
        RECT 94.915 112.905 95.245 113.235 ;
        RECT 106.740 101.420 108.740 211.570 ;
        RECT 112.395 155.065 112.725 155.395 ;
        RECT 112.410 139.075 112.710 155.065 ;
        RECT 112.395 138.745 112.725 139.075 ;
        RECT 106.730 99.570 108.740 101.420 ;
        RECT 121.740 99.720 123.740 211.570 ;
        RECT 121.740 99.570 123.830 99.720 ;
        RECT 31.770 98.150 33.770 99.570 ;
        RECT 9.390 96.150 33.770 98.150 ;
        RECT 9.465 96.095 11.375 96.150 ;
        RECT 106.730 94.060 108.730 99.570 ;
        RECT 121.810 97.750 123.830 99.570 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 6.000 93.980 108.730 94.060 ;
        RECT 6.000 92.060 135.580 93.980 ;
        RECT 106.730 91.980 135.580 92.060 ;
        RECT 106.730 91.960 108.730 91.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

