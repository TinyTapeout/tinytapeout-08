VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_charge_pump
  CLASS BLOCK ;
  FOREIGN tt_um_urish_charge_pump ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.804199 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 22.890999 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 142.200 5.000 143.700 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 151.500 220.100 153.910 223.200 ;
        RECT 151.500 216.410 153.910 219.510 ;
      LAYER nwell ;
        RECT 154.000 215.810 156.410 223.190 ;
      LAYER pwell ;
        RECT 105.900 212.420 110.680 213.320 ;
        RECT 105.900 209.440 106.800 212.420 ;
      LAYER nwell ;
        RECT 106.800 209.440 109.780 212.420 ;
      LAYER pwell ;
        RECT 109.780 209.440 110.680 212.420 ;
        RECT 105.900 208.540 110.680 209.440 ;
        RECT 105.940 184.310 110.720 185.210 ;
        RECT 105.940 181.330 106.840 184.310 ;
      LAYER nwell ;
        RECT 106.840 181.330 109.820 184.310 ;
      LAYER pwell ;
        RECT 109.820 181.330 110.720 184.310 ;
        RECT 105.940 180.430 110.720 181.330 ;
        RECT 105.910 157.270 110.690 158.170 ;
        RECT 105.910 154.290 106.810 157.270 ;
      LAYER nwell ;
        RECT 106.810 154.290 109.790 157.270 ;
      LAYER pwell ;
        RECT 109.790 154.290 110.690 157.270 ;
        RECT 105.910 153.390 110.690 154.290 ;
        RECT 105.910 140.850 110.690 141.750 ;
        RECT 105.910 137.870 106.810 140.850 ;
      LAYER nwell ;
        RECT 106.810 137.870 109.790 140.850 ;
      LAYER pwell ;
        RECT 109.790 137.870 110.690 140.850 ;
        RECT 105.910 136.970 110.690 137.870 ;
      LAYER nwell ;
        RECT 116.000 12.480 158.580 15.870 ;
        RECT 116.000 7.000 158.580 10.390 ;
      LAYER li1 ;
        RECT 151.680 222.850 153.730 223.020 ;
        RECT 151.680 220.450 151.850 222.850 ;
        RECT 152.480 222.340 152.930 222.510 ;
        RECT 152.250 221.130 152.420 222.170 ;
        RECT 152.990 221.130 153.160 222.170 ;
        RECT 152.480 220.790 152.930 220.960 ;
        RECT 153.560 220.450 153.730 222.850 ;
        RECT 151.680 220.280 153.730 220.450 ;
        RECT 154.180 222.840 156.230 223.010 ;
        RECT 154.180 219.850 154.350 222.840 ;
        RECT 154.980 222.330 155.430 222.500 ;
        RECT 154.750 220.575 154.920 222.115 ;
        RECT 155.490 220.575 155.660 222.115 ;
        RECT 154.980 220.190 155.430 220.360 ;
        RECT 156.060 219.850 156.230 222.840 ;
        RECT 154.180 219.680 156.230 219.850 ;
        RECT 151.680 219.160 153.730 219.330 ;
        RECT 151.680 216.760 151.850 219.160 ;
        RECT 152.480 218.650 152.930 218.820 ;
        RECT 152.250 217.440 152.420 218.480 ;
        RECT 152.990 217.440 153.160 218.480 ;
        RECT 152.480 217.100 152.930 217.270 ;
        RECT 153.560 216.760 153.730 219.160 ;
        RECT 151.680 216.590 153.730 216.760 ;
        RECT 154.180 219.150 156.230 219.320 ;
        RECT 154.180 216.160 154.350 219.150 ;
        RECT 154.980 218.640 155.430 218.810 ;
        RECT 154.750 216.885 154.920 218.425 ;
        RECT 155.490 216.885 155.660 218.425 ;
        RECT 154.980 216.500 155.430 216.670 ;
        RECT 156.060 216.160 156.230 219.150 ;
        RECT 154.180 215.990 156.230 216.160 ;
        RECT 106.140 213.020 110.440 213.080 ;
        RECT 105.920 212.910 110.440 213.020 ;
        RECT 105.920 208.950 106.610 212.910 ;
        RECT 107.190 211.860 109.390 212.030 ;
        RECT 107.190 210.000 107.360 211.860 ;
        RECT 107.770 210.490 108.810 211.370 ;
        RECT 109.220 211.360 109.390 211.860 ;
        RECT 109.180 210.620 109.420 211.360 ;
        RECT 109.220 210.000 109.390 210.620 ;
        RECT 107.190 209.830 109.390 210.000 ;
        RECT 110.270 208.950 110.440 212.910 ;
        RECT 105.920 208.900 110.440 208.950 ;
        RECT 106.140 208.780 110.440 208.900 ;
        RECT 106.180 184.900 110.480 184.970 ;
        RECT 105.920 184.800 110.480 184.900 ;
        RECT 105.920 180.840 106.610 184.800 ;
        RECT 107.230 183.750 109.430 183.920 ;
        RECT 107.230 181.890 107.400 183.750 ;
        RECT 109.260 183.280 109.430 183.750 ;
        RECT 107.810 182.380 108.850 183.260 ;
        RECT 109.210 182.420 109.520 183.280 ;
        RECT 109.260 181.890 109.430 182.420 ;
        RECT 107.230 181.720 109.430 181.890 ;
        RECT 110.310 180.840 110.480 184.800 ;
        RECT 105.920 180.780 110.480 180.840 ;
        RECT 106.180 180.670 110.480 180.780 ;
        RECT 106.150 157.840 110.450 157.930 ;
        RECT 105.940 157.760 110.450 157.840 ;
        RECT 105.940 153.800 106.630 157.760 ;
        RECT 107.200 156.710 109.400 156.880 ;
        RECT 107.200 154.850 107.370 156.710 ;
        RECT 109.230 156.300 109.400 156.710 ;
        RECT 107.780 155.340 108.820 156.220 ;
        RECT 109.220 155.410 109.420 156.300 ;
        RECT 109.230 154.850 109.400 155.410 ;
        RECT 107.200 154.680 109.400 154.850 ;
        RECT 110.280 153.800 110.450 157.760 ;
        RECT 105.940 153.720 110.450 153.800 ;
        RECT 106.150 153.630 110.450 153.720 ;
        RECT 106.580 141.510 110.040 141.710 ;
        RECT 106.150 141.340 110.450 141.510 ;
        RECT 106.150 137.380 106.320 141.340 ;
        RECT 106.580 141.240 110.040 141.340 ;
        RECT 107.120 140.290 109.400 140.460 ;
        RECT 107.120 138.430 107.420 140.290 ;
        RECT 107.780 138.920 108.820 139.800 ;
        RECT 109.230 138.430 109.400 140.290 ;
        RECT 107.120 138.320 109.400 138.430 ;
        RECT 107.200 138.260 109.400 138.320 ;
        RECT 110.280 137.380 110.450 141.340 ;
        RECT 106.150 137.210 110.450 137.380 ;
        RECT 116.390 15.310 158.190 15.480 ;
        RECT 116.390 14.740 116.560 15.310 ;
        RECT 116.380 14.510 116.560 14.740 ;
        RECT 117.290 14.620 157.290 14.790 ;
        RECT 116.390 13.040 116.560 14.510 ;
        RECT 117.060 13.945 117.230 14.405 ;
        RECT 157.350 13.945 157.520 14.405 ;
        RECT 117.290 13.560 157.290 13.730 ;
        RECT 158.020 13.040 158.190 15.310 ;
        RECT 116.390 12.870 158.190 13.040 ;
        RECT 116.390 9.830 158.190 10.000 ;
        RECT 116.390 7.560 116.560 9.830 ;
        RECT 117.290 9.140 157.290 9.310 ;
        RECT 117.060 8.465 117.230 8.925 ;
        RECT 157.350 8.465 157.520 8.925 ;
        RECT 117.290 8.080 157.290 8.250 ;
        RECT 158.020 7.560 158.190 9.830 ;
        RECT 116.390 7.390 158.190 7.560 ;
      LAYER met1 ;
        RECT 152.500 222.530 155.400 222.600 ;
        RECT 152.500 222.300 155.410 222.530 ;
        RECT 151.650 221.700 151.880 221.760 ;
        RECT 152.220 221.700 152.450 222.150 ;
        RECT 152.960 221.800 153.190 222.150 ;
        RECT 154.720 221.800 154.950 222.095 ;
        RECT 155.460 221.800 155.690 222.095 ;
        RECT 156.000 221.800 156.300 222.600 ;
        RECT 145.750 221.400 152.450 221.700 ;
        RECT 152.900 221.500 155.000 221.800 ;
        RECT 155.460 221.500 156.300 221.800 ;
        RECT 151.650 221.340 151.880 221.400 ;
        RECT 152.220 221.150 152.450 221.400 ;
        RECT 152.960 221.150 153.190 221.500 ;
        RECT 152.500 220.760 152.910 220.990 ;
        RECT 153.800 219.900 154.100 221.500 ;
        RECT 154.720 220.595 154.950 221.500 ;
        RECT 155.460 220.595 155.690 221.500 ;
        RECT 155.000 220.160 155.410 220.390 ;
        RECT 153.750 219.600 154.150 219.900 ;
        RECT 153.800 218.900 154.100 219.600 ;
        RECT 152.400 218.600 155.500 218.900 ;
        RECT 151.650 218.400 151.880 218.460 ;
        RECT 152.220 218.400 152.450 218.460 ;
        RECT 145.750 218.100 152.450 218.400 ;
        RECT 151.650 218.040 151.880 218.100 ;
        RECT 152.220 217.460 152.450 218.100 ;
        RECT 152.960 218.000 153.190 218.460 ;
        RECT 154.720 218.000 154.950 218.405 ;
        RECT 152.960 217.700 154.950 218.000 ;
        RECT 152.960 217.460 153.190 217.700 ;
        RECT 152.500 217.070 152.910 217.300 ;
        RECT 153.400 215.700 153.700 217.700 ;
        RECT 154.720 216.905 154.950 217.700 ;
        RECT 155.460 218.000 155.690 218.405 ;
        RECT 156.000 218.000 156.300 221.500 ;
        RECT 155.460 217.700 156.300 218.000 ;
        RECT 155.460 216.905 155.690 217.700 ;
        RECT 156.000 217.000 156.300 217.700 ;
        RECT 155.000 216.470 155.410 216.700 ;
        RECT 155.950 216.400 156.350 217.000 ;
        RECT 153.250 214.800 153.950 215.700 ;
        RECT 105.890 213.020 106.640 213.080 ;
        RECT 105.870 208.900 106.660 213.020 ;
        RECT 107.790 210.460 108.790 211.400 ;
        RECT 109.150 211.370 109.450 211.420 ;
        RECT 110.830 211.370 112.550 211.500 ;
        RECT 109.150 210.600 112.550 211.370 ;
        RECT 109.150 210.560 109.450 210.600 ;
        RECT 105.890 208.840 106.640 208.900 ;
        RECT 105.890 184.900 106.640 184.960 ;
        RECT 105.870 180.780 106.660 184.900 ;
        RECT 109.180 183.300 109.550 183.340 ;
        RECT 107.830 183.280 108.830 183.290 ;
        RECT 107.830 182.380 108.840 183.280 ;
        RECT 109.180 182.400 112.550 183.300 ;
        RECT 107.830 182.350 108.830 182.380 ;
        RECT 109.180 182.360 109.550 182.400 ;
        RECT 105.890 180.720 106.640 180.780 ;
        RECT 105.910 157.840 106.660 157.900 ;
        RECT 105.890 153.720 106.680 157.840 ;
        RECT 109.190 156.300 109.450 156.360 ;
        RECT 107.800 155.310 108.800 156.250 ;
        RECT 109.190 155.400 112.570 156.300 ;
        RECT 109.190 155.350 109.450 155.400 ;
        RECT 105.910 153.660 106.660 153.720 ;
        RECT 105.720 141.770 110.640 141.780 ;
        RECT 105.710 141.130 110.640 141.770 ;
        RECT 105.720 141.060 110.640 141.130 ;
        RECT 96.900 140.730 101.100 141.000 ;
        RECT 96.900 140.700 107.480 140.730 ;
        RECT 96.850 139.500 107.480 140.700 ;
        RECT 96.900 138.300 107.480 139.500 ;
        RECT 107.790 138.930 108.800 139.830 ;
        RECT 107.800 138.890 108.800 138.930 ;
        RECT 96.850 138.050 107.480 138.300 ;
        RECT 96.850 137.100 101.100 138.050 ;
        RECT 96.900 135.900 101.100 137.100 ;
        RECT 96.850 134.700 101.100 135.900 ;
        RECT 96.900 134.400 101.100 134.700 ;
        RECT 115.300 14.740 115.680 14.800 ;
        RECT 116.350 14.740 116.590 14.800 ;
        RECT 115.300 14.510 117.145 14.740 ;
        RECT 117.310 14.590 157.270 14.820 ;
        RECT 115.300 14.490 115.680 14.510 ;
        RECT 116.350 14.450 116.590 14.510 ;
        RECT 116.915 14.385 117.145 14.510 ;
        RECT 157.450 14.385 157.650 14.510 ;
        RECT 116.915 13.965 117.260 14.385 ;
        RECT 157.320 13.965 157.650 14.385 ;
        RECT 157.450 13.760 157.650 13.965 ;
        RECT 117.310 13.530 157.650 13.760 ;
        RECT 157.450 11.960 157.650 13.530 ;
        RECT 157.300 11.230 157.740 11.960 ;
        RECT 157.450 10.030 157.650 11.230 ;
        RECT 157.390 9.800 157.710 10.030 ;
        RECT 117.310 9.320 157.270 9.340 ;
        RECT 116.970 9.110 157.270 9.320 ;
        RECT 116.970 8.280 117.480 9.110 ;
        RECT 157.450 8.905 157.650 9.800 ;
        RECT 157.320 8.485 157.650 8.905 ;
        RECT 116.970 8.050 157.270 8.280 ;
        RECT 116.970 5.660 117.480 8.050 ;
        RECT 157.450 7.590 157.650 8.485 ;
        RECT 157.390 7.360 157.710 7.590 ;
        RECT 116.970 5.160 117.490 5.660 ;
        RECT 116.970 5.100 117.480 5.160 ;
      LAYER met2 ;
        RECT 143.750 224.660 144.250 225.260 ;
        RECT 143.850 224.410 144.150 224.660 ;
        RECT 143.850 224.110 154.100 224.410 ;
        RECT 153.800 222.250 154.100 224.110 ;
        RECT 145.800 221.350 146.700 221.750 ;
        RECT 139.500 219.900 140.100 219.950 ;
        RECT 153.800 219.900 154.100 219.950 ;
        RECT 139.500 219.300 154.200 219.900 ;
        RECT 139.500 219.250 140.100 219.300 ;
        RECT 145.800 218.050 146.700 218.450 ;
        RECT 21.600 217.710 25.800 217.990 ;
        RECT 21.040 217.430 25.800 217.710 ;
        RECT 20.480 217.150 25.800 217.430 ;
        RECT 19.920 216.870 25.800 217.150 ;
        RECT 19.640 216.590 25.800 216.870 ;
        RECT 19.360 216.310 25.800 216.590 ;
        RECT 28.600 216.310 31.400 217.430 ;
        RECT 19.080 216.030 25.800 216.310 ;
        RECT 18.800 215.470 25.800 216.030 ;
        RECT 18.520 214.910 25.800 215.470 ;
        RECT 18.240 214.630 25.800 214.910 ;
        RECT 28.880 214.630 31.680 216.310 ;
        RECT 18.240 214.350 22.440 214.630 ;
        RECT 17.960 214.070 21.600 214.350 ;
        RECT 17.960 213.790 21.320 214.070 ;
        RECT 17.960 213.510 21.040 213.790 ;
        RECT 17.960 212.950 20.760 213.510 ;
        RECT 17.960 211.550 20.480 212.950 ;
        RECT 17.960 210.710 20.760 211.550 ;
        RECT 17.960 210.430 21.040 210.710 ;
        RECT 18.240 210.150 21.320 210.430 ;
        RECT 18.240 209.870 21.600 210.150 ;
        RECT 18.240 209.590 22.160 209.870 ;
        RECT 23.280 209.590 25.800 214.630 ;
        RECT 29.160 212.110 31.960 214.630 ;
        RECT 28.880 211.270 31.960 212.110 ;
        RECT 28.600 210.710 31.960 211.270 ;
        RECT 28.320 210.430 31.680 210.710 ;
        RECT 28.040 210.150 31.680 210.430 ;
        RECT 27.760 209.870 31.680 210.150 ;
        RECT 27.200 209.590 31.680 209.870 ;
        RECT 18.520 209.310 25.800 209.590 ;
        RECT 26.640 209.310 31.400 209.590 ;
        RECT 18.520 209.030 31.400 209.310 ;
        RECT 18.800 208.470 31.120 209.030 ;
        RECT 105.920 208.850 106.610 213.070 ;
        RECT 107.850 210.470 108.700 211.420 ;
        RECT 19.080 208.190 30.840 208.470 ;
        RECT 19.360 207.910 30.560 208.190 ;
        RECT 19.640 207.630 30.280 207.910 ;
        RECT 19.920 207.350 30.280 207.630 ;
        RECT 20.200 207.070 29.720 207.350 ;
        RECT 20.760 206.790 29.440 207.070 ;
        RECT 21.320 206.510 28.880 206.790 ;
        RECT 21.880 206.230 28.320 206.510 ;
        RECT 23.000 205.950 27.480 206.230 ;
        RECT 18.240 202.030 20.760 203.990 ;
        RECT 31.960 203.710 33.080 203.990 ;
        RECT 31.120 203.430 34.200 203.710 ;
        RECT 30.560 203.150 34.760 203.430 ;
        RECT 30.280 202.870 35.040 203.150 ;
        RECT 30.000 202.590 35.320 202.870 ;
        RECT 21.600 202.310 23.560 202.590 ;
        RECT 29.720 202.310 35.600 202.590 ;
        RECT 21.040 202.030 24.680 202.310 ;
        RECT 29.720 202.030 35.880 202.310 ;
        RECT 18.240 201.750 25.240 202.030 ;
        RECT 29.440 201.750 35.880 202.030 ;
        RECT 18.240 201.470 25.520 201.750 ;
        RECT 29.440 201.470 36.160 201.750 ;
        RECT 18.240 201.190 25.800 201.470 ;
        RECT 18.240 200.910 26.080 201.190 ;
        RECT 18.240 200.350 26.360 200.910 ;
        RECT 29.160 200.630 36.440 201.470 ;
        RECT 29.160 200.350 36.720 200.630 ;
        RECT 18.240 199.790 26.640 200.350 ;
        RECT 28.880 200.070 32.520 200.350 ;
        RECT 33.360 200.070 36.720 200.350 ;
        RECT 18.240 199.230 26.920 199.790 ;
        RECT 17.960 198.950 21.600 199.230 ;
        RECT 23.560 198.950 26.920 199.230 ;
        RECT 28.880 199.510 31.960 200.070 ;
        RECT 33.640 199.790 36.720 200.070 ;
        RECT 33.920 199.510 37.000 199.790 ;
        RECT 17.960 198.670 21.040 198.950 ;
        RECT 24.120 198.670 27.200 198.950 ;
        RECT 17.960 198.110 20.760 198.670 ;
        RECT 24.400 198.110 27.200 198.670 ;
        RECT 17.960 196.150 20.480 198.110 ;
        RECT 24.680 196.150 27.200 198.110 ;
        RECT 17.960 195.590 20.760 196.150 ;
        RECT 24.400 195.590 27.200 196.150 ;
        RECT 28.880 198.110 31.680 199.510 ;
        RECT 34.200 198.950 37.000 199.510 ;
        RECT 28.880 195.590 31.400 198.110 ;
        RECT 34.480 197.550 37.000 198.950 ;
        RECT 34.760 196.710 37.000 197.550 ;
        RECT 17.960 195.310 21.040 195.590 ;
        RECT 24.120 195.310 26.920 195.590 ;
        RECT 18.240 195.030 21.600 195.310 ;
        RECT 23.560 195.030 26.920 195.310 ;
        RECT 28.600 195.310 31.680 195.590 ;
        RECT 34.480 195.310 37.000 196.710 ;
        RECT 28.600 195.030 31.960 195.310 ;
        RECT 18.240 194.750 27.200 195.030 ;
        RECT 28.320 194.750 31.960 195.030 ;
        RECT 34.200 194.750 37.000 195.310 ;
        RECT 18.240 194.470 27.480 194.750 ;
        RECT 27.760 194.470 32.520 194.750 ;
        RECT 33.920 194.470 37.000 194.750 ;
        RECT 18.520 194.190 37.000 194.470 ;
        RECT 18.520 193.910 36.720 194.190 ;
        RECT 18.800 193.350 36.720 193.910 ;
        RECT 19.080 193.070 36.440 193.350 ;
        RECT 19.360 192.790 36.440 193.070 ;
        RECT 19.640 192.510 36.440 192.790 ;
        RECT 20.200 192.230 24.960 192.510 ;
        RECT 26.080 192.230 30.560 192.510 ;
        RECT 30.840 192.230 36.160 192.510 ;
        RECT 20.480 191.950 24.680 192.230 ;
        RECT 26.360 191.950 30.280 192.230 ;
        RECT 21.600 191.670 23.840 191.950 ;
        RECT 26.920 191.670 29.720 191.950 ;
        RECT 31.120 191.670 35.880 192.230 ;
        RECT 27.760 191.390 29.160 191.670 ;
        RECT 31.680 191.390 35.600 191.670 ;
        RECT 31.960 191.110 35.040 191.390 ;
        RECT 32.520 190.830 34.480 191.110 ;
        RECT 21.040 188.030 31.680 188.310 ;
        RECT 20.200 187.750 31.680 188.030 ;
        RECT 19.640 187.470 31.680 187.750 ;
        RECT 19.360 187.190 31.680 187.470 ;
        RECT 19.080 186.910 31.680 187.190 ;
        RECT 18.800 186.630 31.680 186.910 ;
        RECT 111.600 186.720 112.500 211.550 ;
        RECT 18.520 186.070 31.680 186.630 ;
        RECT 18.240 185.230 31.680 186.070 ;
        RECT 107.810 185.820 112.500 186.720 ;
        RECT 18.240 184.950 30.280 185.230 ;
        RECT 17.960 184.670 22.160 184.950 ;
        RECT 17.960 184.390 21.320 184.670 ;
        RECT 17.960 183.830 21.040 184.390 ;
        RECT 17.960 183.270 20.760 183.830 ;
        RECT 17.960 181.030 20.480 183.270 ;
        RECT 23.280 181.870 25.800 184.950 ;
        RECT 27.480 184.670 30.560 184.950 ;
        RECT 27.760 184.390 30.840 184.670 ;
        RECT 28.040 183.830 31.120 184.390 ;
        RECT 28.320 183.550 31.400 183.830 ;
        RECT 28.600 183.270 31.400 183.550 ;
        RECT 28.880 182.710 31.680 183.270 ;
        RECT 29.160 182.150 31.680 182.710 ;
        RECT 23.280 181.310 26.080 181.870 ;
        RECT 29.160 181.310 31.960 182.150 ;
        RECT 23.280 181.030 26.360 181.310 ;
        RECT 17.960 179.910 20.760 181.030 ;
        RECT 23.560 180.750 26.360 181.030 ;
        RECT 28.880 180.750 31.960 181.310 ;
        RECT 23.560 180.470 26.640 180.750 ;
        RECT 28.600 180.470 31.960 180.750 ;
        RECT 105.920 180.730 106.610 184.950 ;
        RECT 107.810 183.330 108.710 185.820 ;
        RECT 107.810 182.370 108.790 183.330 ;
        RECT 107.890 182.330 108.790 182.370 ;
        RECT 23.560 180.190 27.200 180.470 ;
        RECT 28.040 180.190 31.960 180.470 ;
        RECT 23.560 179.910 31.960 180.190 ;
        RECT 18.240 179.630 20.760 179.910 ;
        RECT 23.840 179.630 31.960 179.910 ;
        RECT 18.240 178.790 21.040 179.630 ;
        RECT 23.840 179.070 31.680 179.630 ;
        RECT 24.120 178.790 31.680 179.070 ;
        RECT 18.520 178.230 21.320 178.790 ;
        RECT 24.120 178.510 31.400 178.790 ;
        RECT 24.400 178.230 31.400 178.510 ;
        RECT 18.520 177.950 21.600 178.230 ;
        RECT 24.680 177.950 31.120 178.230 ;
        RECT 18.800 177.670 21.600 177.950 ;
        RECT 24.960 177.670 30.840 177.950 ;
        RECT 25.240 177.390 30.560 177.670 ;
        RECT 25.520 177.110 30.280 177.390 ;
        RECT 26.080 176.830 29.720 177.110 ;
        RECT 26.920 176.550 28.320 176.830 ;
        RECT 18.240 168.430 20.760 173.470 ;
        RECT 28.600 173.190 31.680 173.470 ;
        RECT 28.880 171.790 31.680 173.190 ;
        RECT 29.160 169.830 31.960 171.790 ;
        RECT 28.880 169.270 31.960 169.830 ;
        RECT 28.600 168.990 31.960 169.270 ;
        RECT 28.320 168.710 31.960 168.990 ;
        RECT 27.760 168.430 31.960 168.710 ;
        RECT 14.040 167.310 31.680 168.430 ;
        RECT 14.040 167.030 31.400 167.310 ;
        RECT 14.320 166.750 31.400 167.030 ;
        RECT 14.320 166.190 31.120 166.750 ;
        RECT 14.600 165.910 30.840 166.190 ;
        RECT 14.600 165.630 30.560 165.910 ;
        RECT 14.600 165.350 30.000 165.630 ;
        RECT 14.600 165.070 29.440 165.350 ;
        RECT 14.880 164.790 27.760 165.070 ;
        RECT 18.240 161.430 20.760 164.790 ;
        RECT 111.600 160.660 112.500 183.350 ;
        RECT 107.810 159.760 112.500 160.660 ;
        RECT 28.880 155.550 31.680 159.470 ;
        RECT 12.920 151.910 31.680 155.550 ;
        RECT 105.940 153.670 106.630 157.890 ;
        RECT 107.810 155.360 108.710 159.760 ;
        RECT 147.900 159.550 148.500 219.300 ;
        RECT 156.000 216.350 156.300 217.050 ;
        RECT 153.300 214.750 153.900 215.750 ;
        RECT 107.850 155.320 108.710 155.360 ;
        RECT 12.920 148.270 15.720 151.910 ;
        RECT 28.880 147.710 31.680 151.910 ;
        RECT 22.440 144.910 26.920 145.190 ;
        RECT 21.600 144.630 28.040 144.910 ;
        RECT 111.680 144.900 112.580 156.280 ;
        RECT 21.040 144.350 28.600 144.630 ;
        RECT 20.480 144.070 29.160 144.350 ;
        RECT 19.920 143.790 29.440 144.070 ;
        RECT 107.840 144.000 112.580 144.900 ;
        RECT 19.640 143.510 30.000 143.790 ;
        RECT 19.360 143.230 30.280 143.510 ;
        RECT 19.080 142.950 30.560 143.230 ;
        RECT 18.800 142.670 30.560 142.950 ;
        RECT 18.800 142.390 30.840 142.670 ;
        RECT 18.520 141.830 31.120 142.390 ;
        RECT 18.240 141.550 31.400 141.830 ;
        RECT 18.240 141.270 23.000 141.550 ;
        RECT 26.640 141.270 31.400 141.550 ;
        RECT 18.240 140.990 22.160 141.270 ;
        RECT 27.480 140.990 31.680 141.270 ;
        RECT 105.760 141.080 106.680 141.820 ;
        RECT 17.960 140.710 21.880 140.990 ;
        RECT 27.760 140.710 31.680 140.990 ;
        RECT 17.960 140.430 21.600 140.710 ;
        RECT 17.960 140.150 21.320 140.430 ;
        RECT 28.320 140.150 31.680 140.710 ;
        RECT 17.960 139.030 21.040 140.150 ;
        RECT 28.600 139.870 31.960 140.150 ;
        RECT 17.960 138.470 20.760 139.030 ;
        RECT 17.960 137.630 21.040 138.470 ;
        RECT 28.880 137.910 31.960 139.870 ;
        RECT 96.900 139.450 98.100 140.750 ;
        RECT 107.840 138.880 108.740 144.000 ;
        RECT 17.960 137.070 21.320 137.630 ;
        RECT 28.600 137.350 31.960 137.910 ;
        RECT 28.320 137.070 31.960 137.350 ;
        RECT 17.960 136.790 21.600 137.070 ;
        RECT 28.320 136.790 31.680 137.070 ;
        RECT 96.900 137.050 98.100 138.350 ;
        RECT 18.240 136.510 21.880 136.790 ;
        RECT 28.040 136.510 31.680 136.790 ;
        RECT 18.240 136.230 22.440 136.510 ;
        RECT 27.480 136.230 31.680 136.510 ;
        RECT 18.240 135.950 23.000 136.230 ;
        RECT 26.920 135.950 31.680 136.230 ;
        RECT 18.520 135.670 24.680 135.950 ;
        RECT 25.240 135.670 31.400 135.950 ;
        RECT 18.520 135.390 31.400 135.670 ;
        RECT 18.800 134.830 31.120 135.390 ;
        RECT 19.080 134.550 30.840 134.830 ;
        RECT 96.900 134.650 98.100 135.950 ;
        RECT 19.360 134.270 30.840 134.550 ;
        RECT 19.640 133.990 30.560 134.270 ;
        RECT 19.920 133.710 30.280 133.990 ;
        RECT 20.200 133.430 30.000 133.710 ;
        RECT 20.760 133.150 29.440 133.430 ;
        RECT 21.040 132.870 28.880 133.150 ;
        RECT 21.880 132.590 28.320 132.870 ;
        RECT 22.720 132.310 27.480 132.590 ;
        RECT 14.320 131.190 15.440 131.470 ;
        RECT 14.320 130.910 16.280 131.190 ;
        RECT 14.320 130.630 17.120 130.910 ;
        RECT 14.320 130.350 17.960 130.630 ;
        RECT 14.320 130.070 19.080 130.350 ;
        RECT 14.320 129.790 19.920 130.070 ;
        RECT 14.320 129.510 20.760 129.790 ;
        RECT 14.320 129.230 21.600 129.510 ;
        RECT 14.320 128.950 22.720 129.230 ;
        RECT 14.320 128.670 23.560 128.950 ;
        RECT 14.320 128.390 24.400 128.670 ;
        RECT 14.320 128.110 25.240 128.390 ;
        RECT 14.320 127.830 26.360 128.110 ;
        RECT 14.880 127.550 27.200 127.830 ;
        RECT 16.000 127.270 28.040 127.550 ;
        RECT 16.840 126.990 29.160 127.270 ;
        RECT 17.960 126.710 30.000 126.990 ;
        RECT 19.080 126.430 30.840 126.710 ;
        RECT 19.920 126.150 31.680 126.430 ;
        RECT 21.040 125.870 31.680 126.150 ;
        RECT 21.880 125.590 31.680 125.870 ;
        RECT 23.000 125.310 31.680 125.590 ;
        RECT 23.840 125.030 31.680 125.310 ;
        RECT 24.960 124.750 31.680 125.030 ;
        RECT 25.800 124.470 31.680 124.750 ;
        RECT 26.920 123.910 31.680 124.470 ;
        RECT 26.080 123.630 31.680 123.910 ;
        RECT 24.960 123.350 31.680 123.630 ;
        RECT 23.840 123.070 31.680 123.350 ;
        RECT 23.000 122.790 31.680 123.070 ;
        RECT 21.880 122.510 31.680 122.790 ;
        RECT 21.040 122.230 31.680 122.510 ;
        RECT 19.920 121.950 31.680 122.230 ;
        RECT 18.800 121.670 31.680 121.950 ;
        RECT 17.960 121.390 30.560 121.670 ;
        RECT 16.840 121.110 29.720 121.390 ;
        RECT 16.000 120.830 28.880 121.110 ;
        RECT 14.880 120.550 28.040 120.830 ;
        RECT 14.320 120.270 26.920 120.550 ;
        RECT 14.320 119.990 26.080 120.270 ;
        RECT 14.320 119.710 25.240 119.990 ;
        RECT 14.320 119.430 24.400 119.710 ;
        RECT 14.320 119.150 23.280 119.430 ;
        RECT 14.320 118.870 22.440 119.150 ;
        RECT 14.320 118.590 21.600 118.870 ;
        RECT 14.320 118.310 20.480 118.590 ;
        RECT 14.320 118.030 19.640 118.310 ;
        RECT 14.320 117.750 18.800 118.030 ;
        RECT 14.320 117.470 17.960 117.750 ;
        RECT 14.320 117.190 16.840 117.470 ;
        RECT 14.320 116.910 16.000 117.190 ;
        RECT 14.320 116.630 15.160 116.910 ;
        RECT 20.760 100.110 31.680 100.390 ;
        RECT 19.920 99.830 31.680 100.110 ;
        RECT 19.360 99.550 31.680 99.830 ;
        RECT 19.080 99.270 31.680 99.550 ;
        RECT 18.800 98.990 31.680 99.270 ;
        RECT 18.520 98.430 31.680 98.990 ;
        RECT 18.240 97.870 31.680 98.430 ;
        RECT 17.960 97.030 31.680 97.870 ;
        RECT 17.960 96.750 21.880 97.030 ;
        RECT 17.960 96.470 21.320 96.750 ;
        RECT 17.960 95.910 21.040 96.470 ;
        RECT 17.960 95.350 20.760 95.910 ;
        RECT 17.960 94.510 21.040 95.350 ;
        RECT 18.240 94.230 21.320 94.510 ;
        RECT 18.240 93.950 21.600 94.230 ;
        RECT 18.520 93.670 21.880 93.950 ;
        RECT 18.520 93.390 22.160 93.670 ;
        RECT 18.800 93.110 22.440 93.390 ;
        RECT 19.080 92.830 22.720 93.110 ;
        RECT 19.360 92.550 23.000 92.830 ;
        RECT 12.920 89.190 31.680 92.550 ;
        RECT 18.240 84.990 20.760 86.670 ;
        RECT 31.400 86.390 33.640 86.670 ;
        RECT 30.840 86.110 34.480 86.390 ;
        RECT 30.280 85.830 34.760 86.110 ;
        RECT 30.000 85.550 35.040 85.830 ;
        RECT 30.000 85.270 35.320 85.550 ;
        RECT 21.320 84.990 24.120 85.270 ;
        RECT 29.720 84.990 35.600 85.270 ;
        RECT 18.240 84.710 24.960 84.990 ;
        RECT 29.440 84.710 35.880 84.990 ;
        RECT 18.240 84.430 25.240 84.710 ;
        RECT 18.240 84.150 25.520 84.430 ;
        RECT 29.440 84.150 36.160 84.710 ;
        RECT 18.240 83.870 25.800 84.150 ;
        RECT 18.240 83.590 26.080 83.870 ;
        RECT 29.160 83.590 36.440 84.150 ;
        RECT 18.240 83.310 26.360 83.590 ;
        RECT 29.160 83.310 36.720 83.590 ;
        RECT 18.240 82.750 26.640 83.310 ;
        RECT 28.880 83.030 36.720 83.310 ;
        RECT 28.880 82.750 32.240 83.030 ;
        RECT 33.360 82.750 36.720 83.030 ;
        RECT 18.240 82.190 26.920 82.750 ;
        RECT 18.240 81.910 22.160 82.190 ;
        RECT 23.000 81.910 26.920 82.190 ;
        RECT 17.960 81.630 21.320 81.910 ;
        RECT 23.840 81.630 26.920 81.910 ;
        RECT 28.880 82.470 31.960 82.750 ;
        RECT 33.920 82.470 36.720 82.750 ;
        RECT 17.960 81.350 21.040 81.630 ;
        RECT 24.120 81.350 27.200 81.630 ;
        RECT 17.960 81.070 20.760 81.350 ;
        RECT 24.400 81.070 27.200 81.350 ;
        RECT 17.960 78.830 20.480 81.070 ;
        RECT 24.680 78.830 27.200 81.070 ;
        RECT 17.960 78.550 20.760 78.830 ;
        RECT 17.960 78.270 21.040 78.550 ;
        RECT 24.400 78.270 27.200 78.830 ;
        RECT 28.880 81.070 31.680 82.470 ;
        RECT 34.200 81.630 37.000 82.470 ;
        RECT 28.880 78.550 31.400 81.070 ;
        RECT 34.480 80.230 37.000 81.630 ;
        RECT 34.760 79.670 37.000 80.230 ;
        RECT 28.600 78.270 31.400 78.550 ;
        RECT 34.480 78.270 37.000 79.670 ;
        RECT 17.960 77.990 21.320 78.270 ;
        RECT 23.840 77.990 26.920 78.270 ;
        RECT 28.600 77.990 31.680 78.270 ;
        RECT 18.240 77.710 21.880 77.990 ;
        RECT 23.280 77.710 26.920 77.990 ;
        RECT 28.320 77.710 31.960 77.990 ;
        RECT 34.200 77.710 37.000 78.270 ;
        RECT 18.240 77.430 27.200 77.710 ;
        RECT 28.320 77.430 32.240 77.710 ;
        RECT 33.920 77.430 37.000 77.710 ;
        RECT 18.240 77.150 32.800 77.430 ;
        RECT 33.640 77.150 37.000 77.430 ;
        RECT 18.520 76.590 36.720 77.150 ;
        RECT 18.800 76.310 36.720 76.590 ;
        RECT 19.080 76.030 36.720 76.310 ;
        RECT 19.080 75.750 36.440 76.030 ;
        RECT 19.360 75.470 36.440 75.750 ;
        RECT 19.920 75.190 25.240 75.470 ;
        RECT 25.800 75.190 36.160 75.470 ;
        RECT 20.200 74.910 24.960 75.190 ;
        RECT 26.080 74.910 30.280 75.190 ;
        RECT 30.840 74.910 36.160 75.190 ;
        RECT 20.760 74.630 24.400 74.910 ;
        RECT 26.640 74.630 30.000 74.910 ;
        RECT 31.120 74.630 35.880 74.910 ;
        RECT 27.200 74.350 29.440 74.630 ;
        RECT 31.400 74.350 35.600 74.630 ;
        RECT 31.680 74.070 35.320 74.350 ;
        RECT 32.240 73.790 34.760 74.070 ;
        RECT 13.760 67.630 15.440 67.910 ;
        RECT 28.880 67.630 31.680 71.550 ;
        RECT 13.200 67.350 16.000 67.630 ;
        RECT 12.920 67.070 16.280 67.350 ;
        RECT 12.640 66.510 16.560 67.070 ;
        RECT 12.640 66.230 16.840 66.510 ;
        RECT 12.360 65.110 16.840 66.230 ;
        RECT 12.640 64.830 16.840 65.110 ;
        RECT 12.640 64.270 16.560 64.830 ;
        RECT 12.920 63.990 16.280 64.270 ;
        RECT 18.240 63.990 31.680 67.630 ;
        RECT 13.200 63.710 16.000 63.990 ;
        RECT 13.760 63.430 15.440 63.710 ;
        RECT 18.240 60.350 20.760 63.990 ;
        RECT 28.880 59.790 31.680 63.990 ;
        RECT 14.320 53.630 31.680 56.990 ;
        RECT 21.320 48.030 24.120 53.630 ;
        RECT 14.320 44.670 31.680 48.030 ;
        RECT 35.880 39.070 37.000 39.350 ;
        RECT 35.320 38.790 37.560 39.070 ;
        RECT 34.760 38.510 37.840 38.790 ;
        RECT 34.480 38.230 37.840 38.510 ;
        RECT 33.920 37.950 37.840 38.230 ;
        RECT 33.360 37.670 37.840 37.950 ;
        RECT 32.800 37.390 37.840 37.670 ;
        RECT 32.520 37.110 37.840 37.390 ;
        RECT 31.960 36.830 37.840 37.110 ;
        RECT 31.400 36.550 37.840 36.830 ;
        RECT 31.120 36.270 37.840 36.550 ;
        RECT 30.560 35.990 37.840 36.270 ;
        RECT 30.000 35.710 37.840 35.990 ;
        RECT 29.440 35.430 37.840 35.710 ;
        RECT 29.160 35.150 37.840 35.430 ;
        RECT 28.600 34.870 34.480 35.150 ;
        RECT 28.040 34.590 34.200 34.870 ;
        RECT 27.480 34.310 33.640 34.590 ;
        RECT 27.200 34.030 33.080 34.310 ;
        RECT 26.640 33.750 32.520 34.030 ;
        RECT 26.080 33.470 32.240 33.750 ;
        RECT 25.520 33.190 31.680 33.470 ;
        RECT 25.240 32.910 31.120 33.190 ;
        RECT 24.680 32.630 30.840 32.910 ;
        RECT 24.120 32.350 30.280 32.630 ;
        RECT 23.840 32.070 29.720 32.350 ;
        RECT 23.280 31.790 29.160 32.070 ;
        RECT 22.720 31.510 28.880 31.790 ;
        RECT 22.160 31.230 28.320 31.510 ;
        RECT 21.880 30.950 27.760 31.230 ;
        RECT 21.320 30.670 27.200 30.950 ;
        RECT 20.760 30.390 26.920 30.670 ;
        RECT 20.200 30.110 26.360 30.390 ;
        RECT 19.920 29.830 25.800 30.110 ;
        RECT 19.360 29.550 25.240 29.830 ;
        RECT 18.800 29.270 24.960 29.550 ;
        RECT 18.240 28.990 24.400 29.270 ;
        RECT 17.960 28.710 23.840 28.990 ;
        RECT 17.400 28.430 23.560 28.710 ;
        RECT 16.840 28.150 23.000 28.430 ;
        RECT 16.560 27.870 22.440 28.150 ;
        RECT 16.000 27.590 21.880 27.870 ;
        RECT 15.440 27.310 21.600 27.590 ;
        RECT 14.880 27.030 21.040 27.310 ;
        RECT 14.600 26.750 20.480 27.030 ;
        RECT 14.040 26.470 19.920 26.750 ;
        RECT 13.480 26.190 19.640 26.470 ;
        RECT 12.920 25.910 19.080 26.190 ;
        RECT 12.640 25.630 18.520 25.910 ;
        RECT 23.000 25.630 23.560 25.910 ;
        RECT 12.080 25.350 17.960 25.630 ;
        RECT 23.000 25.350 24.400 25.630 ;
        RECT 11.520 25.070 17.680 25.350 ;
        RECT 23.280 25.070 25.520 25.350 ;
        RECT 10.960 24.790 17.120 25.070 ;
        RECT 23.280 24.790 26.640 25.070 ;
        RECT 10.680 24.510 16.560 24.790 ;
        RECT 23.560 24.510 27.480 24.790 ;
        RECT 30.560 24.510 31.120 24.790 ;
        RECT 10.120 24.230 16.280 24.510 ;
        RECT 17.960 24.230 18.800 24.510 ;
        RECT 23.560 24.230 28.600 24.510 ;
        RECT 30.840 24.230 31.680 24.510 ;
        RECT 9.560 23.950 15.720 24.230 ;
        RECT 17.960 23.950 19.360 24.230 ;
        RECT 23.840 23.950 29.440 24.230 ;
        RECT 30.840 23.950 31.960 24.230 ;
        RECT 9.280 23.670 15.160 23.950 ;
        RECT 17.960 23.670 20.200 23.950 ;
        RECT 23.840 23.670 30.560 23.950 ;
        RECT 31.120 23.670 32.520 23.950 ;
        RECT 9.000 23.390 14.600 23.670 ;
        RECT 17.960 23.390 20.760 23.670 ;
        RECT 24.120 23.390 32.800 23.670 ;
        RECT 9.000 23.110 14.320 23.390 ;
        RECT 17.960 23.110 21.600 23.390 ;
        RECT 24.120 23.110 33.360 23.390 ;
        RECT 9.000 22.830 13.760 23.110 ;
        RECT 17.960 22.830 22.440 23.110 ;
        RECT 24.400 22.830 33.640 23.110 ;
        RECT 9.000 22.550 13.480 22.830 ;
        RECT 17.960 22.550 23.000 22.830 ;
        RECT 24.400 22.550 26.080 22.830 ;
        RECT 26.920 22.550 34.200 22.830 ;
        RECT 9.000 22.270 14.040 22.550 ;
        RECT 17.960 22.270 23.840 22.550 ;
        RECT 24.680 22.270 26.360 22.550 ;
        RECT 28.320 22.270 34.480 22.550 ;
        RECT 9.000 21.990 14.320 22.270 ;
        RECT 9.000 21.710 14.880 21.990 ;
        RECT 17.960 21.710 26.360 22.270 ;
        RECT 30.000 21.990 34.760 22.270 ;
        RECT 30.560 21.710 34.480 21.990 ;
        RECT 9.280 21.430 15.440 21.710 ;
        RECT 9.840 21.150 15.720 21.430 ;
        RECT 17.960 21.150 26.640 21.710 ;
        RECT 30.280 21.430 33.080 21.710 ;
        RECT 30.000 21.150 31.680 21.430 ;
        RECT 10.400 20.870 16.280 21.150 ;
        RECT 19.080 20.870 26.920 21.150 ;
        RECT 30.000 20.870 30.560 21.150 ;
        RECT 10.680 20.590 16.840 20.870 ;
        RECT 19.920 20.590 26.920 20.870 ;
        RECT 11.240 20.310 17.400 20.590 ;
        RECT 21.040 20.310 27.200 20.590 ;
        RECT 11.800 20.030 17.680 20.310 ;
        RECT 21.880 20.030 27.200 20.310 ;
        RECT 12.360 19.750 18.240 20.030 ;
        RECT 23.000 19.750 27.480 20.030 ;
        RECT 12.640 19.470 18.800 19.750 ;
        RECT 24.120 19.470 27.480 19.750 ;
        RECT 13.200 19.190 19.360 19.470 ;
        RECT 24.960 19.190 27.760 19.470 ;
        RECT 13.760 18.910 19.640 19.190 ;
        RECT 26.080 18.910 27.760 19.190 ;
        RECT 14.320 18.630 20.200 18.910 ;
        RECT 27.200 18.630 27.760 18.910 ;
        RECT 14.600 18.350 20.760 18.630 ;
        RECT 15.160 18.070 21.320 18.350 ;
        RECT 15.720 17.790 21.600 18.070 ;
        RECT 16.000 17.510 22.160 17.790 ;
        RECT 16.560 17.230 22.720 17.510 ;
        RECT 17.120 16.950 23.000 17.230 ;
        RECT 17.680 16.670 23.560 16.950 ;
        RECT 17.960 16.390 24.120 16.670 ;
        RECT 18.520 16.110 24.680 16.390 ;
        RECT 19.080 15.830 24.960 16.110 ;
        RECT 19.640 15.550 25.520 15.830 ;
        RECT 19.920 15.270 26.080 15.550 ;
        RECT 20.480 14.990 26.640 15.270 ;
        RECT 21.040 14.710 26.920 14.990 ;
        RECT 21.600 14.430 27.480 14.710 ;
        RECT 21.880 14.150 28.040 14.430 ;
        RECT 22.440 13.870 28.600 14.150 ;
        RECT 23.000 13.590 28.880 13.870 ;
        RECT 23.280 13.310 29.440 13.590 ;
        RECT 23.840 13.030 30.000 13.310 ;
        RECT 24.400 12.750 30.280 13.030 ;
        RECT 24.960 12.470 30.840 12.750 ;
        RECT 25.240 12.190 31.400 12.470 ;
        RECT 25.800 11.910 31.960 12.190 ;
        RECT 26.360 11.630 32.240 11.910 ;
        RECT 26.920 11.350 32.800 11.630 ;
        RECT 27.200 11.070 33.360 11.350 ;
        RECT 27.760 10.790 33.920 11.070 ;
        RECT 28.320 10.510 34.200 10.790 ;
        RECT 28.880 10.230 34.760 10.510 ;
        RECT 35.040 10.230 37.840 35.150 ;
        RECT 115.350 14.440 115.630 14.850 ;
        RECT 157.350 11.180 157.690 12.010 ;
        RECT 29.160 9.950 37.840 10.230 ;
        RECT 29.720 9.670 37.840 9.950 ;
        RECT 30.280 9.390 37.840 9.670 ;
        RECT 30.560 9.110 37.840 9.390 ;
        RECT 31.120 8.830 37.840 9.110 ;
        RECT 31.680 8.550 37.840 8.830 ;
        RECT 32.240 8.270 37.840 8.550 ;
        RECT 32.520 7.990 37.840 8.270 ;
        RECT 33.080 7.710 37.840 7.990 ;
        RECT 33.640 7.430 37.840 7.710 ;
        RECT 34.200 7.150 37.840 7.430 ;
        RECT 34.480 6.870 37.840 7.150 ;
        RECT 35.040 6.590 37.840 6.870 ;
        RECT 35.600 6.310 37.280 6.590 ;
        RECT 49.500 5.700 50.100 5.750 ;
        RECT 117.020 5.700 117.440 5.710 ;
        RECT 49.500 5.100 117.470 5.700 ;
        RECT 49.500 5.050 50.100 5.100 ;
      LAYER met3 ;
        RECT 143.700 224.685 144.300 225.235 ;
        RECT 145.450 222.500 147.050 223.500 ;
        RECT 139.450 219.275 140.150 219.925 ;
        RECT 107.800 217.500 143.200 218.400 ;
        RECT 145.500 218.000 147.000 222.500 ;
        RECT 105.870 208.875 106.660 213.045 ;
        RECT 107.800 211.395 108.700 217.500 ;
        RECT 142.300 217.200 143.200 217.500 ;
        RECT 142.160 217.000 143.750 217.200 ;
        RECT 155.950 217.000 156.350 217.025 ;
        RECT 142.160 216.400 156.350 217.000 ;
        RECT 142.160 216.300 143.750 216.400 ;
        RECT 155.950 216.375 156.350 216.400 ;
        RECT 142.300 216.230 143.200 216.300 ;
        RECT 107.800 210.495 108.750 211.395 ;
        RECT 111.550 210.575 112.550 211.525 ;
        RECT 107.800 210.440 108.700 210.495 ;
        RECT 113.500 189.500 139.995 215.500 ;
        RECT 153.250 214.775 153.950 215.725 ;
        RECT 105.870 180.755 106.660 184.925 ;
        RECT 111.550 182.375 112.550 183.325 ;
        RECT 113.400 162.300 139.895 188.300 ;
        RECT 153.300 187.200 153.900 214.775 ;
        RECT 140.350 186.600 153.900 187.200 ;
        RECT 105.890 153.695 106.680 157.865 ;
        RECT 111.760 155.455 112.540 156.235 ;
        RECT 64.200 119.700 95.695 145.700 ;
        RECT 105.710 141.105 106.730 141.795 ;
        RECT 96.900 140.725 98.100 141.000 ;
        RECT 96.850 139.475 98.150 140.725 ;
        RECT 96.900 138.325 98.100 139.475 ;
        RECT 96.850 137.075 98.150 138.325 ;
        RECT 96.900 135.925 98.100 137.075 ;
        RECT 96.850 134.675 98.150 135.925 ;
        RECT 113.400 135.000 139.895 161.000 ;
        RECT 147.850 160.200 148.550 160.225 ;
        RECT 140.350 159.600 148.550 160.200 ;
        RECT 147.850 159.575 148.550 159.600 ;
        RECT 96.900 15.680 98.100 134.675 ;
        RECT 96.900 14.825 115.650 15.680 ;
        RECT 96.900 14.480 115.680 14.825 ;
        RECT 115.300 14.465 115.680 14.480 ;
        RECT 157.300 11.205 157.740 11.985 ;
        RECT 49.450 5.075 50.150 5.725 ;
      LAYER met4 ;
        RECT 143.745 224.760 143.830 225.215 ;
        RECT 144.130 224.760 144.255 225.215 ;
        RECT 30.670 223.500 30.970 224.760 ;
        RECT 33.430 223.500 33.730 224.760 ;
        RECT 36.190 223.500 36.490 224.760 ;
        RECT 38.950 223.500 39.250 224.760 ;
        RECT 41.710 223.500 42.010 224.760 ;
        RECT 44.470 223.500 44.770 224.760 ;
        RECT 47.230 223.500 47.530 224.760 ;
        RECT 49.990 223.500 50.290 224.760 ;
        RECT 52.750 223.500 53.050 224.760 ;
        RECT 55.510 223.500 55.810 224.760 ;
        RECT 58.270 223.500 58.570 224.760 ;
        RECT 61.030 223.500 61.330 224.760 ;
        RECT 63.790 223.500 64.090 224.760 ;
        RECT 66.550 223.500 66.850 224.760 ;
        RECT 69.310 223.500 69.610 224.760 ;
        RECT 72.070 223.500 72.370 224.760 ;
        RECT 74.830 223.500 75.130 224.760 ;
        RECT 77.590 223.500 77.890 224.760 ;
        RECT 80.350 223.500 80.650 224.760 ;
        RECT 83.110 223.500 83.410 224.760 ;
        RECT 85.870 223.500 86.170 224.760 ;
        RECT 88.630 223.500 88.930 224.760 ;
        RECT 91.390 223.500 91.690 224.760 ;
        RECT 94.150 223.500 94.450 224.760 ;
        RECT 143.745 224.705 144.255 224.760 ;
        RECT 145.495 223.500 147.005 223.505 ;
        RECT 30.630 222.500 147.005 223.500 ;
        RECT 49.000 220.760 50.500 222.500 ;
        RECT 64.895 139.200 94.505 145.005 ;
        RECT 95.195 141.000 95.675 145.640 ;
        RECT 105.730 141.080 106.730 222.500 ;
        RECT 145.495 222.495 147.005 222.500 ;
        RECT 139.495 219.295 140.105 219.905 ;
        RECT 139.500 215.440 140.100 219.295 ;
        RECT 142.195 216.295 142.200 217.205 ;
        RECT 143.700 216.295 143.705 217.205 ;
        RECT 139.495 215.100 140.100 215.440 ;
        RECT 111.595 211.500 112.505 211.505 ;
        RECT 114.195 211.500 138.805 214.805 ;
        RECT 111.595 210.600 138.805 211.500 ;
        RECT 111.595 210.595 112.505 210.600 ;
        RECT 114.195 190.195 138.805 210.600 ;
        RECT 139.495 189.560 139.975 215.100 ;
        RECT 139.395 188.100 139.875 188.240 ;
        RECT 111.595 183.300 112.505 183.305 ;
        RECT 114.095 183.300 138.705 187.605 ;
        RECT 111.595 182.400 138.705 183.300 ;
        RECT 111.595 182.395 112.505 182.400 ;
        RECT 114.095 162.995 138.705 182.400 ;
        RECT 139.395 186.000 141.600 188.100 ;
        RECT 139.395 162.360 139.875 186.000 ;
        RECT 139.395 160.800 139.875 160.940 ;
        RECT 114.095 156.300 138.705 160.305 ;
        RECT 111.760 155.400 138.705 156.300 ;
        RECT 50.500 128.400 94.505 139.200 ;
        RECT 95.100 140.705 98.100 141.000 ;
        RECT 95.100 139.495 98.105 140.705 ;
        RECT 95.100 138.305 98.100 139.495 ;
        RECT 95.100 137.095 98.105 138.305 ;
        RECT 95.100 135.905 98.100 137.095 ;
        RECT 95.100 134.695 98.105 135.905 ;
        RECT 114.095 135.695 138.705 155.400 ;
        RECT 139.395 159.000 141.600 160.800 ;
        RECT 139.395 135.060 139.875 159.000 ;
        RECT 95.100 134.400 98.100 134.695 ;
        RECT 64.895 120.395 94.505 128.400 ;
        RECT 95.195 119.760 95.675 134.400 ;
        RECT 156.410 11.140 157.770 12.040 ;
        RECT 156.410 3.900 157.310 11.140 ;
        RECT 151.810 3.000 157.310 3.900 ;
        RECT 151.810 1.000 152.710 3.000 ;
  END
END tt_um_urish_charge_pump
END LIBRARY

