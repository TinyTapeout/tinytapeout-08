module tt_um_tommythorn_maxbw (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input VPWR;
 input VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire net145;
 wire \tokenflow_inst.i1.c.q ;
 wire \tokenflow_inst.i10.cg.b ;
 wire \tokenflow_inst.i10.cg.q ;
 wire \tokenflow_inst.i10.d0.inv_chain[0] ;
 wire \tokenflow_inst.i10.d0.inv_chain[1] ;
 wire \tokenflow_inst.i11.i.cg.q ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[0] ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[1] ;
 wire \tokenflow_inst.i2.cg1.q ;
 wire \tokenflow_inst.i2.cg2.a ;
 wire \tokenflow_inst.i2.cg2.q ;
 wire \tokenflow_inst.i2.cg3.q ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i3.ydata[0] ;
 wire \tokenflow_inst.i3.ydata[10] ;
 wire \tokenflow_inst.i3.ydata[11] ;
 wire \tokenflow_inst.i3.ydata[12] ;
 wire \tokenflow_inst.i3.ydata[13] ;
 wire \tokenflow_inst.i3.ydata[14] ;
 wire \tokenflow_inst.i3.ydata[15] ;
 wire \tokenflow_inst.i3.ydata[16] ;
 wire \tokenflow_inst.i3.ydata[17] ;
 wire \tokenflow_inst.i3.ydata[18] ;
 wire \tokenflow_inst.i3.ydata[19] ;
 wire \tokenflow_inst.i3.ydata[1] ;
 wire \tokenflow_inst.i3.ydata[20] ;
 wire \tokenflow_inst.i3.ydata[21] ;
 wire \tokenflow_inst.i3.ydata[22] ;
 wire \tokenflow_inst.i3.ydata[23] ;
 wire \tokenflow_inst.i3.ydata[24] ;
 wire \tokenflow_inst.i3.ydata[25] ;
 wire \tokenflow_inst.i3.ydata[26] ;
 wire \tokenflow_inst.i3.ydata[27] ;
 wire \tokenflow_inst.i3.ydata[28] ;
 wire \tokenflow_inst.i3.ydata[29] ;
 wire \tokenflow_inst.i3.ydata[2] ;
 wire \tokenflow_inst.i3.ydata[30] ;
 wire \tokenflow_inst.i3.ydata[31] ;
 wire \tokenflow_inst.i3.ydata[32] ;
 wire \tokenflow_inst.i3.ydata[33] ;
 wire \tokenflow_inst.i3.ydata[34] ;
 wire \tokenflow_inst.i3.ydata[35] ;
 wire \tokenflow_inst.i3.ydata[36] ;
 wire \tokenflow_inst.i3.ydata[37] ;
 wire \tokenflow_inst.i3.ydata[38] ;
 wire \tokenflow_inst.i3.ydata[39] ;
 wire \tokenflow_inst.i3.ydata[3] ;
 wire \tokenflow_inst.i3.ydata[40] ;
 wire \tokenflow_inst.i3.ydata[41] ;
 wire \tokenflow_inst.i3.ydata[42] ;
 wire \tokenflow_inst.i3.ydata[43] ;
 wire \tokenflow_inst.i3.ydata[44] ;
 wire \tokenflow_inst.i3.ydata[45] ;
 wire \tokenflow_inst.i3.ydata[46] ;
 wire \tokenflow_inst.i3.ydata[47] ;
 wire \tokenflow_inst.i3.ydata[48] ;
 wire \tokenflow_inst.i3.ydata[49] ;
 wire \tokenflow_inst.i3.ydata[4] ;
 wire \tokenflow_inst.i3.ydata[50] ;
 wire \tokenflow_inst.i3.ydata[51] ;
 wire \tokenflow_inst.i3.ydata[52] ;
 wire \tokenflow_inst.i3.ydata[53] ;
 wire \tokenflow_inst.i3.ydata[54] ;
 wire \tokenflow_inst.i3.ydata[55] ;
 wire \tokenflow_inst.i3.ydata[56] ;
 wire \tokenflow_inst.i3.ydata[57] ;
 wire \tokenflow_inst.i3.ydata[58] ;
 wire \tokenflow_inst.i3.ydata[59] ;
 wire \tokenflow_inst.i3.ydata[5] ;
 wire \tokenflow_inst.i3.ydata[60] ;
 wire \tokenflow_inst.i3.ydata[61] ;
 wire \tokenflow_inst.i3.ydata[62] ;
 wire \tokenflow_inst.i3.ydata[63] ;
 wire \tokenflow_inst.i3.ydata[64] ;
 wire \tokenflow_inst.i3.ydata[65] ;
 wire \tokenflow_inst.i3.ydata[66] ;
 wire \tokenflow_inst.i3.ydata[67] ;
 wire \tokenflow_inst.i3.ydata[68] ;
 wire \tokenflow_inst.i3.ydata[69] ;
 wire \tokenflow_inst.i3.ydata[6] ;
 wire \tokenflow_inst.i3.ydata[70] ;
 wire \tokenflow_inst.i3.ydata[71] ;
 wire \tokenflow_inst.i3.ydata[72] ;
 wire \tokenflow_inst.i3.ydata[73] ;
 wire \tokenflow_inst.i3.ydata[74] ;
 wire \tokenflow_inst.i3.ydata[75] ;
 wire \tokenflow_inst.i3.ydata[76] ;
 wire \tokenflow_inst.i3.ydata[77] ;
 wire \tokenflow_inst.i3.ydata[7] ;
 wire \tokenflow_inst.i3.ydata[8] ;
 wire \tokenflow_inst.i3.ydata[9] ;
 wire \tokenflow_inst.i6.cg_elem.q ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i6.ydata[0] ;
 wire \tokenflow_inst.i6.ydata[10] ;
 wire \tokenflow_inst.i6.ydata[11] ;
 wire \tokenflow_inst.i6.ydata[12] ;
 wire \tokenflow_inst.i6.ydata[13] ;
 wire \tokenflow_inst.i6.ydata[14] ;
 wire \tokenflow_inst.i6.ydata[15] ;
 wire \tokenflow_inst.i6.ydata[16] ;
 wire \tokenflow_inst.i6.ydata[17] ;
 wire \tokenflow_inst.i6.ydata[18] ;
 wire \tokenflow_inst.i6.ydata[19] ;
 wire \tokenflow_inst.i6.ydata[1] ;
 wire \tokenflow_inst.i6.ydata[20] ;
 wire \tokenflow_inst.i6.ydata[21] ;
 wire \tokenflow_inst.i6.ydata[22] ;
 wire \tokenflow_inst.i6.ydata[23] ;
 wire \tokenflow_inst.i6.ydata[24] ;
 wire \tokenflow_inst.i6.ydata[25] ;
 wire \tokenflow_inst.i6.ydata[26] ;
 wire \tokenflow_inst.i6.ydata[27] ;
 wire \tokenflow_inst.i6.ydata[28] ;
 wire \tokenflow_inst.i6.ydata[29] ;
 wire \tokenflow_inst.i6.ydata[2] ;
 wire \tokenflow_inst.i6.ydata[30] ;
 wire \tokenflow_inst.i6.ydata[31] ;
 wire \tokenflow_inst.i6.ydata[32] ;
 wire \tokenflow_inst.i6.ydata[33] ;
 wire \tokenflow_inst.i6.ydata[34] ;
 wire \tokenflow_inst.i6.ydata[35] ;
 wire \tokenflow_inst.i6.ydata[36] ;
 wire \tokenflow_inst.i6.ydata[37] ;
 wire \tokenflow_inst.i6.ydata[38] ;
 wire \tokenflow_inst.i6.ydata[39] ;
 wire \tokenflow_inst.i6.ydata[3] ;
 wire \tokenflow_inst.i6.ydata[40] ;
 wire \tokenflow_inst.i6.ydata[41] ;
 wire \tokenflow_inst.i6.ydata[42] ;
 wire \tokenflow_inst.i6.ydata[43] ;
 wire \tokenflow_inst.i6.ydata[44] ;
 wire \tokenflow_inst.i6.ydata[45] ;
 wire \tokenflow_inst.i6.ydata[46] ;
 wire \tokenflow_inst.i6.ydata[47] ;
 wire \tokenflow_inst.i6.ydata[48] ;
 wire \tokenflow_inst.i6.ydata[49] ;
 wire \tokenflow_inst.i6.ydata[4] ;
 wire \tokenflow_inst.i6.ydata[50] ;
 wire \tokenflow_inst.i6.ydata[51] ;
 wire \tokenflow_inst.i6.ydata[52] ;
 wire \tokenflow_inst.i6.ydata[53] ;
 wire \tokenflow_inst.i6.ydata[54] ;
 wire \tokenflow_inst.i6.ydata[55] ;
 wire \tokenflow_inst.i6.ydata[56] ;
 wire \tokenflow_inst.i6.ydata[57] ;
 wire \tokenflow_inst.i6.ydata[58] ;
 wire \tokenflow_inst.i6.ydata[59] ;
 wire \tokenflow_inst.i6.ydata[5] ;
 wire \tokenflow_inst.i6.ydata[60] ;
 wire \tokenflow_inst.i6.ydata[61] ;
 wire \tokenflow_inst.i6.ydata[62] ;
 wire \tokenflow_inst.i6.ydata[63] ;
 wire \tokenflow_inst.i6.ydata[64] ;
 wire \tokenflow_inst.i6.ydata[65] ;
 wire \tokenflow_inst.i6.ydata[66] ;
 wire \tokenflow_inst.i6.ydata[67] ;
 wire \tokenflow_inst.i6.ydata[68] ;
 wire \tokenflow_inst.i6.ydata[69] ;
 wire \tokenflow_inst.i6.ydata[6] ;
 wire \tokenflow_inst.i6.ydata[70] ;
 wire \tokenflow_inst.i6.ydata[71] ;
 wire \tokenflow_inst.i6.ydata[72] ;
 wire \tokenflow_inst.i6.ydata[73] ;
 wire \tokenflow_inst.i6.ydata[74] ;
 wire \tokenflow_inst.i6.ydata[75] ;
 wire \tokenflow_inst.i6.ydata[76] ;
 wire \tokenflow_inst.i6.ydata[77] ;
 wire \tokenflow_inst.i6.ydata[7] ;
 wire \tokenflow_inst.i6.ydata[8] ;
 wire \tokenflow_inst.i6.ydata[9] ;
 wire \tokenflow_inst.i78.cg_elem.q ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i78.ydata[0] ;
 wire \tokenflow_inst.i78.ydata[10] ;
 wire \tokenflow_inst.i78.ydata[11] ;
 wire \tokenflow_inst.i78.ydata[12] ;
 wire \tokenflow_inst.i78.ydata[13] ;
 wire \tokenflow_inst.i78.ydata[14] ;
 wire \tokenflow_inst.i78.ydata[15] ;
 wire \tokenflow_inst.i78.ydata[16] ;
 wire \tokenflow_inst.i78.ydata[17] ;
 wire \tokenflow_inst.i78.ydata[18] ;
 wire \tokenflow_inst.i78.ydata[19] ;
 wire \tokenflow_inst.i78.ydata[1] ;
 wire \tokenflow_inst.i78.ydata[20] ;
 wire \tokenflow_inst.i78.ydata[21] ;
 wire \tokenflow_inst.i78.ydata[22] ;
 wire \tokenflow_inst.i78.ydata[23] ;
 wire \tokenflow_inst.i78.ydata[24] ;
 wire \tokenflow_inst.i78.ydata[25] ;
 wire \tokenflow_inst.i78.ydata[26] ;
 wire \tokenflow_inst.i78.ydata[27] ;
 wire \tokenflow_inst.i78.ydata[28] ;
 wire \tokenflow_inst.i78.ydata[29] ;
 wire \tokenflow_inst.i78.ydata[2] ;
 wire \tokenflow_inst.i78.ydata[30] ;
 wire \tokenflow_inst.i78.ydata[31] ;
 wire \tokenflow_inst.i78.ydata[32] ;
 wire \tokenflow_inst.i78.ydata[33] ;
 wire \tokenflow_inst.i78.ydata[34] ;
 wire \tokenflow_inst.i78.ydata[35] ;
 wire \tokenflow_inst.i78.ydata[36] ;
 wire \tokenflow_inst.i78.ydata[37] ;
 wire \tokenflow_inst.i78.ydata[38] ;
 wire \tokenflow_inst.i78.ydata[39] ;
 wire \tokenflow_inst.i78.ydata[3] ;
 wire \tokenflow_inst.i78.ydata[40] ;
 wire \tokenflow_inst.i78.ydata[41] ;
 wire \tokenflow_inst.i78.ydata[42] ;
 wire \tokenflow_inst.i78.ydata[43] ;
 wire \tokenflow_inst.i78.ydata[44] ;
 wire \tokenflow_inst.i78.ydata[45] ;
 wire \tokenflow_inst.i78.ydata[46] ;
 wire \tokenflow_inst.i78.ydata[47] ;
 wire \tokenflow_inst.i78.ydata[48] ;
 wire \tokenflow_inst.i78.ydata[49] ;
 wire \tokenflow_inst.i78.ydata[4] ;
 wire \tokenflow_inst.i78.ydata[50] ;
 wire \tokenflow_inst.i78.ydata[51] ;
 wire \tokenflow_inst.i78.ydata[52] ;
 wire \tokenflow_inst.i78.ydata[53] ;
 wire \tokenflow_inst.i78.ydata[54] ;
 wire \tokenflow_inst.i78.ydata[55] ;
 wire \tokenflow_inst.i78.ydata[56] ;
 wire \tokenflow_inst.i78.ydata[57] ;
 wire \tokenflow_inst.i78.ydata[58] ;
 wire \tokenflow_inst.i78.ydata[59] ;
 wire \tokenflow_inst.i78.ydata[5] ;
 wire \tokenflow_inst.i78.ydata[60] ;
 wire \tokenflow_inst.i78.ydata[61] ;
 wire \tokenflow_inst.i78.ydata[62] ;
 wire \tokenflow_inst.i78.ydata[63] ;
 wire \tokenflow_inst.i78.ydata[64] ;
 wire \tokenflow_inst.i78.ydata[65] ;
 wire \tokenflow_inst.i78.ydata[66] ;
 wire \tokenflow_inst.i78.ydata[67] ;
 wire \tokenflow_inst.i78.ydata[68] ;
 wire \tokenflow_inst.i78.ydata[69] ;
 wire \tokenflow_inst.i78.ydata[6] ;
 wire \tokenflow_inst.i78.ydata[70] ;
 wire \tokenflow_inst.i78.ydata[71] ;
 wire \tokenflow_inst.i78.ydata[72] ;
 wire \tokenflow_inst.i78.ydata[73] ;
 wire \tokenflow_inst.i78.ydata[74] ;
 wire \tokenflow_inst.i78.ydata[75] ;
 wire \tokenflow_inst.i78.ydata[76] ;
 wire \tokenflow_inst.i78.ydata[77] ;
 wire \tokenflow_inst.i78.ydata[7] ;
 wire \tokenflow_inst.i78.ydata[8] ;
 wire \tokenflow_inst.i78.ydata[9] ;
 wire \tokenflow_inst.i8.cg_elem.q ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i8.ydata[0] ;
 wire \tokenflow_inst.i8.ydata[10] ;
 wire \tokenflow_inst.i8.ydata[11] ;
 wire \tokenflow_inst.i8.ydata[12] ;
 wire \tokenflow_inst.i8.ydata[13] ;
 wire \tokenflow_inst.i8.ydata[14] ;
 wire \tokenflow_inst.i8.ydata[15] ;
 wire \tokenflow_inst.i8.ydata[16] ;
 wire \tokenflow_inst.i8.ydata[17] ;
 wire \tokenflow_inst.i8.ydata[18] ;
 wire \tokenflow_inst.i8.ydata[19] ;
 wire \tokenflow_inst.i8.ydata[1] ;
 wire \tokenflow_inst.i8.ydata[20] ;
 wire \tokenflow_inst.i8.ydata[21] ;
 wire \tokenflow_inst.i8.ydata[22] ;
 wire \tokenflow_inst.i8.ydata[23] ;
 wire \tokenflow_inst.i8.ydata[24] ;
 wire \tokenflow_inst.i8.ydata[25] ;
 wire \tokenflow_inst.i8.ydata[26] ;
 wire \tokenflow_inst.i8.ydata[27] ;
 wire \tokenflow_inst.i8.ydata[28] ;
 wire \tokenflow_inst.i8.ydata[29] ;
 wire \tokenflow_inst.i8.ydata[2] ;
 wire \tokenflow_inst.i8.ydata[30] ;
 wire \tokenflow_inst.i8.ydata[31] ;
 wire \tokenflow_inst.i8.ydata[32] ;
 wire \tokenflow_inst.i8.ydata[33] ;
 wire \tokenflow_inst.i8.ydata[34] ;
 wire \tokenflow_inst.i8.ydata[35] ;
 wire \tokenflow_inst.i8.ydata[36] ;
 wire \tokenflow_inst.i8.ydata[37] ;
 wire \tokenflow_inst.i8.ydata[38] ;
 wire \tokenflow_inst.i8.ydata[39] ;
 wire \tokenflow_inst.i8.ydata[3] ;
 wire \tokenflow_inst.i8.ydata[40] ;
 wire \tokenflow_inst.i8.ydata[41] ;
 wire \tokenflow_inst.i8.ydata[42] ;
 wire \tokenflow_inst.i8.ydata[43] ;
 wire \tokenflow_inst.i8.ydata[44] ;
 wire \tokenflow_inst.i8.ydata[45] ;
 wire \tokenflow_inst.i8.ydata[46] ;
 wire \tokenflow_inst.i8.ydata[47] ;
 wire \tokenflow_inst.i8.ydata[48] ;
 wire \tokenflow_inst.i8.ydata[49] ;
 wire \tokenflow_inst.i8.ydata[4] ;
 wire \tokenflow_inst.i8.ydata[50] ;
 wire \tokenflow_inst.i8.ydata[51] ;
 wire \tokenflow_inst.i8.ydata[52] ;
 wire \tokenflow_inst.i8.ydata[53] ;
 wire \tokenflow_inst.i8.ydata[54] ;
 wire \tokenflow_inst.i8.ydata[55] ;
 wire \tokenflow_inst.i8.ydata[56] ;
 wire \tokenflow_inst.i8.ydata[57] ;
 wire \tokenflow_inst.i8.ydata[58] ;
 wire \tokenflow_inst.i8.ydata[59] ;
 wire \tokenflow_inst.i8.ydata[5] ;
 wire \tokenflow_inst.i8.ydata[60] ;
 wire \tokenflow_inst.i8.ydata[61] ;
 wire \tokenflow_inst.i8.ydata[62] ;
 wire \tokenflow_inst.i8.ydata[63] ;
 wire \tokenflow_inst.i8.ydata[64] ;
 wire \tokenflow_inst.i8.ydata[65] ;
 wire \tokenflow_inst.i8.ydata[66] ;
 wire \tokenflow_inst.i8.ydata[67] ;
 wire \tokenflow_inst.i8.ydata[68] ;
 wire \tokenflow_inst.i8.ydata[69] ;
 wire \tokenflow_inst.i8.ydata[6] ;
 wire \tokenflow_inst.i8.ydata[70] ;
 wire \tokenflow_inst.i8.ydata[71] ;
 wire \tokenflow_inst.i8.ydata[72] ;
 wire \tokenflow_inst.i8.ydata[73] ;
 wire \tokenflow_inst.i8.ydata[74] ;
 wire \tokenflow_inst.i8.ydata[75] ;
 wire \tokenflow_inst.i8.ydata[76] ;
 wire \tokenflow_inst.i8.ydata[77] ;
 wire \tokenflow_inst.i8.ydata[7] ;
 wire \tokenflow_inst.i8.ydata[8] ;
 wire \tokenflow_inst.i8.ydata[9] ;
 wire \tokenflow_inst.i9.c.q ;
 wire \tokenflow_inst.ii1.cg_elem.q ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii1.ydata[0] ;
 wire \tokenflow_inst.ii1.ydata[10] ;
 wire \tokenflow_inst.ii1.ydata[11] ;
 wire \tokenflow_inst.ii1.ydata[12] ;
 wire \tokenflow_inst.ii1.ydata[13] ;
 wire \tokenflow_inst.ii1.ydata[14] ;
 wire \tokenflow_inst.ii1.ydata[15] ;
 wire \tokenflow_inst.ii1.ydata[16] ;
 wire \tokenflow_inst.ii1.ydata[17] ;
 wire \tokenflow_inst.ii1.ydata[18] ;
 wire \tokenflow_inst.ii1.ydata[19] ;
 wire \tokenflow_inst.ii1.ydata[1] ;
 wire \tokenflow_inst.ii1.ydata[20] ;
 wire \tokenflow_inst.ii1.ydata[21] ;
 wire \tokenflow_inst.ii1.ydata[22] ;
 wire \tokenflow_inst.ii1.ydata[23] ;
 wire \tokenflow_inst.ii1.ydata[24] ;
 wire \tokenflow_inst.ii1.ydata[25] ;
 wire \tokenflow_inst.ii1.ydata[2] ;
 wire \tokenflow_inst.ii1.ydata[3] ;
 wire \tokenflow_inst.ii1.ydata[4] ;
 wire \tokenflow_inst.ii1.ydata[5] ;
 wire \tokenflow_inst.ii1.ydata[6] ;
 wire \tokenflow_inst.ii1.ydata[7] ;
 wire \tokenflow_inst.ii1.ydata[8] ;
 wire \tokenflow_inst.ii1.ydata[9] ;
 wire \tokenflow_inst.ii2.cg_elem.q ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii2.ydata[0] ;
 wire \tokenflow_inst.ii2.ydata[10] ;
 wire \tokenflow_inst.ii2.ydata[11] ;
 wire \tokenflow_inst.ii2.ydata[12] ;
 wire \tokenflow_inst.ii2.ydata[13] ;
 wire \tokenflow_inst.ii2.ydata[14] ;
 wire \tokenflow_inst.ii2.ydata[15] ;
 wire \tokenflow_inst.ii2.ydata[16] ;
 wire \tokenflow_inst.ii2.ydata[17] ;
 wire \tokenflow_inst.ii2.ydata[18] ;
 wire \tokenflow_inst.ii2.ydata[19] ;
 wire \tokenflow_inst.ii2.ydata[1] ;
 wire \tokenflow_inst.ii2.ydata[20] ;
 wire \tokenflow_inst.ii2.ydata[21] ;
 wire \tokenflow_inst.ii2.ydata[22] ;
 wire \tokenflow_inst.ii2.ydata[23] ;
 wire \tokenflow_inst.ii2.ydata[24] ;
 wire \tokenflow_inst.ii2.ydata[25] ;
 wire \tokenflow_inst.ii2.ydata[2] ;
 wire \tokenflow_inst.ii2.ydata[3] ;
 wire \tokenflow_inst.ii2.ydata[4] ;
 wire \tokenflow_inst.ii2.ydata[5] ;
 wire \tokenflow_inst.ii2.ydata[6] ;
 wire \tokenflow_inst.ii2.ydata[7] ;
 wire \tokenflow_inst.ii2.ydata[8] ;
 wire \tokenflow_inst.ii2.ydata[9] ;
 wire \tokenflow_inst.ii3.i.cg_elem.q ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii3.i.ydata[0] ;
 wire \tokenflow_inst.ii3.i.ydata[10] ;
 wire \tokenflow_inst.ii3.i.ydata[11] ;
 wire \tokenflow_inst.ii3.i.ydata[12] ;
 wire \tokenflow_inst.ii3.i.ydata[13] ;
 wire \tokenflow_inst.ii3.i.ydata[14] ;
 wire \tokenflow_inst.ii3.i.ydata[15] ;
 wire \tokenflow_inst.ii3.i.ydata[16] ;
 wire \tokenflow_inst.ii3.i.ydata[17] ;
 wire \tokenflow_inst.ii3.i.ydata[18] ;
 wire \tokenflow_inst.ii3.i.ydata[19] ;
 wire \tokenflow_inst.ii3.i.ydata[1] ;
 wire \tokenflow_inst.ii3.i.ydata[20] ;
 wire \tokenflow_inst.ii3.i.ydata[21] ;
 wire \tokenflow_inst.ii3.i.ydata[22] ;
 wire \tokenflow_inst.ii3.i.ydata[23] ;
 wire \tokenflow_inst.ii3.i.ydata[24] ;
 wire \tokenflow_inst.ii3.i.ydata[25] ;
 wire \tokenflow_inst.ii3.i.ydata[2] ;
 wire \tokenflow_inst.ii3.i.ydata[3] ;
 wire \tokenflow_inst.ii3.i.ydata[4] ;
 wire \tokenflow_inst.ii3.i.ydata[5] ;
 wire \tokenflow_inst.ii3.i.ydata[6] ;
 wire \tokenflow_inst.ii3.i.ydata[7] ;
 wire \tokenflow_inst.ii3.i.ydata[8] ;
 wire \tokenflow_inst.ii3.i.ydata[9] ;
 wire \tokenflow_inst.ii4.c.q ;
 wire net137;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;

 sky130_fd_sc_hd__inv_2 _0792_ (.A(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _0793_ (.A(net86),
    .B(\tokenflow_inst.i2.cg1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0777_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(\tokenflow_inst.ii3.i.ydata[0] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _0795_ (.A(net118),
    .B(\tokenflow_inst.i2.cg1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0778_));
 sky130_fd_sc_hd__a21o_1 _0796_ (.A1(\tokenflow_inst.i78.ydata[0] ),
    .A2(net9),
    .B1(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _0797_ (.A(\tokenflow_inst.ii3.i.ydata[1] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _0798_ (.A1(\tokenflow_inst.i78.ydata[1] ),
    .A2(net9),
    .B1(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _0799_ (.A1(\tokenflow_inst.ii3.i.ydata[2] ),
    .A2(net19),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_1 _0800_ (.A1(\tokenflow_inst.ii3.i.ydata[3] ),
    .A2(net19),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _0801_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(net20),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _0802_ (.A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(net20),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _0803_ (.A1(\tokenflow_inst.ii3.i.ydata[6] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\tokenflow_inst.ii3.i.ydata[7] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(\tokenflow_inst.ii3.i.ydata[8] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _0806_ (.A1(\tokenflow_inst.ii3.i.ydata[9] ),
    .A2(net16),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(\tokenflow_inst.ii3.i.ydata[11] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(\tokenflow_inst.ii3.i.ydata[12] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _0810_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _0811_ (.A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _0812_ (.A1(\tokenflow_inst.ii3.i.ydata[15] ),
    .A2(net15),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_1 _0813_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(net15),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(\tokenflow_inst.ii3.i.ydata[17] ),
    .A2(net15),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _0816_ (.A1(\tokenflow_inst.ii3.i.ydata[19] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _0818_ (.A1(\tokenflow_inst.ii3.i.ydata[21] ),
    .A2(net15),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(net14),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _0820_ (.A1(\tokenflow_inst.ii3.i.ydata[23] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _0821_ (.A(\tokenflow_inst.ii3.i.ydata[24] ),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__a21o_1 _0822_ (.A1(\tokenflow_inst.i78.ydata[24] ),
    .A2(net5),
    .B1(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _0823_ (.A(\tokenflow_inst.ii3.i.ydata[25] ),
    .B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_1 _0824_ (.A1(\tokenflow_inst.i78.ydata[25] ),
    .A2(net5),
    .B1(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__a21o_1 _0825_ (.A1(\tokenflow_inst.i78.ydata[26] ),
    .A2(net8),
    .B1(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__a21o_1 _0826_ (.A1(\tokenflow_inst.i78.ydata[27] ),
    .A2(net8),
    .B1(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _0827_ (.A1(\tokenflow_inst.ii3.i.ydata[2] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\tokenflow_inst.ii3.i.ydata[3] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _0829_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _0830_ (.A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _0831_ (.A1(\tokenflow_inst.ii3.i.ydata[6] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__a22o_1 _0832_ (.A1(\tokenflow_inst.ii3.i.ydata[7] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(\tokenflow_inst.ii3.i.ydata[8] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0834_ (.A1(\tokenflow_inst.ii3.i.ydata[9] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0835_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _0836_ (.A1(\tokenflow_inst.ii3.i.ydata[11] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_1 _0837_ (.A1(\tokenflow_inst.ii3.i.ydata[12] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _0838_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _0839_ (.A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0840_ (.A1(\tokenflow_inst.ii3.i.ydata[15] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(\tokenflow_inst.ii3.i.ydata[17] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _0843_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(\tokenflow_inst.ii3.i.ydata[19] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_1 _0845_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(net16),
    .B1(net11),
    .B2(\tokenflow_inst.i78.ydata[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _0846_ (.A1(\tokenflow_inst.ii3.i.ydata[21] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_1 _0847_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(net16),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _0848_ (.A1(\tokenflow_inst.ii3.i.ydata[23] ),
    .A2(net13),
    .B1(net4),
    .B2(\tokenflow_inst.i78.ydata[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _0849_ (.A1(\tokenflow_inst.ii3.i.ydata[2] ),
    .A2(net19),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\tokenflow_inst.ii3.i.ydata[3] ),
    .A2(net19),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _0851_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(net20),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(net20),
    .B1(net9),
    .B2(\tokenflow_inst.i78.ydata[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _0853_ (.A1(\tokenflow_inst.ii3.i.ydata[6] ),
    .A2(net18),
    .B1(net8),
    .B2(\tokenflow_inst.i78.ydata[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\tokenflow_inst.ii3.i.ydata[7] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _0855_ (.A1(\tokenflow_inst.ii3.i.ydata[8] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(\tokenflow_inst.ii3.i.ydata[9] ),
    .A2(net17),
    .B1(net7),
    .B2(\tokenflow_inst.i78.ydata[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__a22o_1 _0857_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(net13),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_1 _0858_ (.A1(\tokenflow_inst.ii3.i.ydata[11] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(\tokenflow_inst.ii3.i.ydata[12] ),
    .A2(net12),
    .B1(net3),
    .B2(\tokenflow_inst.i78.ydata[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _0860_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0861_ (.A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_1 _0862_ (.A1(\tokenflow_inst.ii3.i.ydata[15] ),
    .A2(net14),
    .B1(net5),
    .B2(\tokenflow_inst.i78.ydata[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _0863_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(net14),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0864_ (.A1(\tokenflow_inst.ii3.i.ydata[17] ),
    .A2(net14),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _0865_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_1 _0866_ (.A1(\tokenflow_inst.ii3.i.ydata[19] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0867_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(net20),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(\tokenflow_inst.ii3.i.ydata[21] ),
    .A2(net19),
    .B1(net10),
    .B2(\tokenflow_inst.i78.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _0869_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(net15),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _0870_ (.A1(\tokenflow_inst.ii3.i.ydata[23] ),
    .A2(net14),
    .B1(net6),
    .B2(\tokenflow_inst.i78.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__a21o_1 _0871_ (.A1(\tokenflow_inst.i78.ydata[76] ),
    .A2(net5),
    .B1(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(\tokenflow_inst.i78.ydata[77] ),
    .A2(net5),
    .B1(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _0873_ (.A(net118),
    .B(\tokenflow_inst.ii4.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _0874_ (.A(net86),
    .B(\tokenflow_inst.ii2.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0353_));
 sky130_fd_sc_hd__a21o_1 _0875_ (.A1(\tokenflow_inst.ii2.d0_elem.inv_chain[2] ),
    .A2(\tokenflow_inst.ii2.cg_elem.q ),
    .B1(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _0876_ (.A(net116),
    .B(\tokenflow_inst.ii2.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(net116),
    .B(\tokenflow_inst.ii2.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _0878_ (.A(net118),
    .B(\tokenflow_inst.ii2.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(net118),
    .B(\tokenflow_inst.ii2.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__and2_1 _0880_ (.A(net117),
    .B(\tokenflow_inst.ii2.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__and2_1 _0881_ (.A(net117),
    .B(\tokenflow_inst.ii2.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _0882_ (.A(net145),
    .B(\tokenflow_inst.ii2.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__and2_1 _0883_ (.A(net114),
    .B(\tokenflow_inst.ii2.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _0884_ (.A(net111),
    .B(\tokenflow_inst.ii2.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(net114),
    .B(\tokenflow_inst.ii2.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _0886_ (.A(net90),
    .B(\tokenflow_inst.ii2.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(net92),
    .B(\tokenflow_inst.ii2.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _0888_ (.A(net95),
    .B(\tokenflow_inst.ii2.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _0889_ (.A(net95),
    .B(\tokenflow_inst.ii2.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(net95),
    .B(\tokenflow_inst.ii2.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(net94),
    .B(\tokenflow_inst.ii2.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _0892_ (.A(net99),
    .B(\tokenflow_inst.ii2.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__and2_1 _0893_ (.A(net97),
    .B(\tokenflow_inst.ii2.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _0894_ (.A(net110),
    .B(\tokenflow_inst.ii2.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(net110),
    .B(\tokenflow_inst.ii2.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _0896_ (.A(net113),
    .B(\tokenflow_inst.ii2.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _0897_ (.A(net113),
    .B(\tokenflow_inst.ii2.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__and2_1 _0898_ (.A(net99),
    .B(\tokenflow_inst.ii2.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _0899_ (.A(net99),
    .B(\tokenflow_inst.ii2.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _0900_ (.A(net99),
    .B(\tokenflow_inst.ii2.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _0901_ (.A(net94),
    .B(\tokenflow_inst.ii2.ydata[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__and2_1 _0902_ (.A(net116),
    .B(\tokenflow_inst.ii1.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _0903_ (.A(net116),
    .B(\tokenflow_inst.ii1.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(net118),
    .B(\tokenflow_inst.ii1.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _0905_ (.A(net118),
    .B(\tokenflow_inst.ii1.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__and2_1 _0906_ (.A(net117),
    .B(\tokenflow_inst.ii1.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__and2_1 _0907_ (.A(net117),
    .B(\tokenflow_inst.ii1.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _0908_ (.A(net111),
    .B(\tokenflow_inst.ii1.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(net114),
    .B(\tokenflow_inst.ii1.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _0910_ (.A(net111),
    .B(\tokenflow_inst.ii1.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(net113),
    .B(\tokenflow_inst.ii1.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _0912_ (.A(net91),
    .B(\tokenflow_inst.ii1.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _0913_ (.A(net92),
    .B(\tokenflow_inst.ii1.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _0914_ (.A(net95),
    .B(\tokenflow_inst.ii1.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__and2_1 _0915_ (.A(net95),
    .B(\tokenflow_inst.ii1.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _0916_ (.A(net95),
    .B(\tokenflow_inst.ii1.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(net94),
    .B(\tokenflow_inst.ii1.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _0918_ (.A(net100),
    .B(\tokenflow_inst.ii1.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _0919_ (.A(net97),
    .B(\tokenflow_inst.ii1.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _0920_ (.A(net110),
    .B(\tokenflow_inst.ii1.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(net112),
    .B(\tokenflow_inst.ii1.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _0922_ (.A(net113),
    .B(\tokenflow_inst.ii1.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(net113),
    .B(\tokenflow_inst.ii1.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _0924_ (.A(net99),
    .B(\tokenflow_inst.ii1.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _0925_ (.A(net94),
    .B(\tokenflow_inst.ii1.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _0926_ (.A(net94),
    .B(\tokenflow_inst.ii1.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _0927_ (.A(net94),
    .B(\tokenflow_inst.ii1.ydata[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _0928_ (.A(net86),
    .B(\tokenflow_inst.ii3.i.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__o21ai_1 _0929_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .B1(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0779_));
 sky130_fd_sc_hd__a21oi_1 _0930_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .B1(_0779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0011_));
 sky130_fd_sc_hd__a21oi_1 _0931_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .B1(\tokenflow_inst.ii3.i.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0780_));
 sky130_fd_sc_hd__a31o_1 _0932_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .A3(\tokenflow_inst.ii3.i.ydata[2] ),
    .B1(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_1 _0933_ (.A(_0780_),
    .B(_0781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0018_));
 sky130_fd_sc_hd__a31o_1 _0934_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .A3(\tokenflow_inst.ii3.i.ydata[2] ),
    .B1(\tokenflow_inst.ii3.i.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0782_));
 sky130_fd_sc_hd__and4_1 _0935_ (.A(\tokenflow_inst.ii3.i.ydata[0] ),
    .B(\tokenflow_inst.ii3.i.ydata[1] ),
    .C(\tokenflow_inst.ii3.i.ydata[2] ),
    .D(\tokenflow_inst.ii3.i.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0783_));
 sky130_fd_sc_hd__and3b_1 _0936_ (.A_N(_0783_),
    .B(net117),
    .C(_0782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__a21oi_1 _0937_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(_0783_),
    .B1(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0784_));
 sky130_fd_sc_hd__o21a_1 _0938_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(_0783_),
    .B1(_0784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__a21o_1 _0939_ (.A1(\tokenflow_inst.ii3.i.ydata[4] ),
    .A2(_0783_),
    .B1(\tokenflow_inst.ii3.i.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0785_));
 sky130_fd_sc_hd__and3_1 _0940_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(\tokenflow_inst.ii3.i.ydata[5] ),
    .C(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0786_));
 sky130_fd_sc_hd__and3b_1 _0941_ (.A_N(_0786_),
    .B(net114),
    .C(_0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__and4_1 _0942_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(\tokenflow_inst.ii3.i.ydata[5] ),
    .C(\tokenflow_inst.ii3.i.ydata[6] ),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_1 _0943_ (.A1(\tokenflow_inst.ii3.i.ydata[6] ),
    .A2(_0786_),
    .B1(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_1 _0944_ (.A(_0787_),
    .B(_0788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0022_));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(\tokenflow_inst.ii3.i.ydata[7] ),
    .B(_0787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0789_));
 sky130_fd_sc_hd__o21ai_1 _0946_ (.A1(\tokenflow_inst.ii3.i.ydata[7] ),
    .A2(_0787_),
    .B1(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _0947_ (.A(_0789_),
    .B(_0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0023_));
 sky130_fd_sc_hd__and3_1 _0948_ (.A(\tokenflow_inst.ii3.i.ydata[7] ),
    .B(\tokenflow_inst.ii3.i.ydata[8] ),
    .C(_0787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0791_));
 sky130_fd_sc_hd__o21ai_1 _0949_ (.A1(\tokenflow_inst.ii3.i.ydata[8] ),
    .A2(_0789_),
    .B1(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0411_));
 sky130_fd_sc_hd__nor2_1 _0950_ (.A(_0791_),
    .B(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0024_));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(\tokenflow_inst.ii3.i.ydata[9] ),
    .B(_0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__and4_2 _0952_ (.A(\tokenflow_inst.ii3.i.ydata[7] ),
    .B(\tokenflow_inst.ii3.i.ydata[8] ),
    .C(\tokenflow_inst.ii3.i.ydata[9] ),
    .D(_0787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__and3b_1 _0953_ (.A_N(_0413_),
    .B(net113),
    .C(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__a21oi_1 _0954_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(_0413_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0414_));
 sky130_fd_sc_hd__o21a_1 _0955_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(_0413_),
    .B1(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__a21o_1 _0956_ (.A1(\tokenflow_inst.ii3.i.ydata[10] ),
    .A2(_0413_),
    .B1(\tokenflow_inst.ii3.i.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__and3_1 _0957_ (.A(\tokenflow_inst.ii3.i.ydata[10] ),
    .B(\tokenflow_inst.ii3.i.ydata[11] ),
    .C(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__and3b_1 _0958_ (.A_N(_0416_),
    .B(net91),
    .C(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__and4_2 _0959_ (.A(\tokenflow_inst.ii3.i.ydata[10] ),
    .B(\tokenflow_inst.ii3.i.ydata[11] ),
    .C(\tokenflow_inst.ii3.i.ydata[12] ),
    .D(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__o21ai_1 _0960_ (.A1(\tokenflow_inst.ii3.i.ydata[12] ),
    .A2(_0416_),
    .B1(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _0961_ (.A(_0417_),
    .B(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0003_));
 sky130_fd_sc_hd__a21oi_1 _0962_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(_0417_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0419_));
 sky130_fd_sc_hd__o21a_1 _0963_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(_0417_),
    .B1(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__a21oi_1 _0964_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(_0417_),
    .B1(\tokenflow_inst.ii3.i.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0420_));
 sky130_fd_sc_hd__a31o_1 _0965_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(\tokenflow_inst.ii3.i.ydata[14] ),
    .A3(_0417_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__nor2_1 _0966_ (.A(_0420_),
    .B(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0005_));
 sky130_fd_sc_hd__a31o_1 _0967_ (.A1(\tokenflow_inst.ii3.i.ydata[13] ),
    .A2(\tokenflow_inst.ii3.i.ydata[14] ),
    .A3(_0417_),
    .B1(\tokenflow_inst.ii3.i.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__and4_2 _0968_ (.A(\tokenflow_inst.ii3.i.ydata[13] ),
    .B(\tokenflow_inst.ii3.i.ydata[14] ),
    .C(\tokenflow_inst.ii3.i.ydata[15] ),
    .D(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__and3b_1 _0969_ (.A_N(_0423_),
    .B(net95),
    .C(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__a21oi_1 _0970_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(_0423_),
    .B1(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0424_));
 sky130_fd_sc_hd__o21a_1 _0971_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(_0423_),
    .B1(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__a21o_1 _0972_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(_0423_),
    .B1(\tokenflow_inst.ii3.i.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__and3_1 _0973_ (.A(\tokenflow_inst.ii3.i.ydata[16] ),
    .B(\tokenflow_inst.ii3.i.ydata[17] ),
    .C(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__and3b_1 _0974_ (.A_N(_0426_),
    .B(net97),
    .C(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__o21ai_1 _0975_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(_0426_),
    .B1(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0427_));
 sky130_fd_sc_hd__a21oi_1 _0976_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(_0426_),
    .B1(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0009_));
 sky130_fd_sc_hd__a21o_1 _0977_ (.A1(\tokenflow_inst.ii3.i.ydata[18] ),
    .A2(_0426_),
    .B1(\tokenflow_inst.ii3.i.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__and2_1 _0978_ (.A(\tokenflow_inst.ii3.i.ydata[18] ),
    .B(\tokenflow_inst.ii3.i.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__and4_1 _0979_ (.A(\tokenflow_inst.ii3.i.ydata[16] ),
    .B(\tokenflow_inst.ii3.i.ydata[17] ),
    .C(_0423_),
    .D(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__and3b_1 _0980_ (.A_N(_0430_),
    .B(net100),
    .C(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _0981_ (.A(\tokenflow_inst.ii3.i.ydata[20] ),
    .B(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__o21ai_1 _0982_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(_0430_),
    .B1(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0432_));
 sky130_fd_sc_hd__nor2_1 _0983_ (.A(_0431_),
    .B(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0012_));
 sky130_fd_sc_hd__and3_1 _0984_ (.A(\tokenflow_inst.ii3.i.ydata[20] ),
    .B(\tokenflow_inst.ii3.i.ydata[21] ),
    .C(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__o21ai_1 _0985_ (.A1(\tokenflow_inst.ii3.i.ydata[21] ),
    .A2(_0431_),
    .B1(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0434_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(_0433_),
    .B(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0013_));
 sky130_fd_sc_hd__and2_1 _0987_ (.A(\tokenflow_inst.ii3.i.ydata[22] ),
    .B(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__o21ai_1 _0988_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(_0433_),
    .B1(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(_0435_),
    .B(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0014_));
 sky130_fd_sc_hd__a21oi_1 _0990_ (.A1(\tokenflow_inst.ii3.i.ydata[23] ),
    .A2(_0435_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0437_));
 sky130_fd_sc_hd__o21a_1 _0991_ (.A1(\tokenflow_inst.ii3.i.ydata[23] ),
    .A2(_0435_),
    .B1(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__a31o_1 _0992_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(\tokenflow_inst.ii3.i.ydata[23] ),
    .A3(_0433_),
    .B1(\tokenflow_inst.ii3.i.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _0993_ (.A(\tokenflow_inst.ii3.i.ydata[23] ),
    .B(\tokenflow_inst.ii3.i.ydata[24] ),
    .C(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__and3b_1 _0994_ (.A_N(_0439_),
    .B(net94),
    .C(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__o21ai_1 _0995_ (.A1(\tokenflow_inst.ii3.i.ydata[25] ),
    .A2(_0439_),
    .B1(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0440_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(\tokenflow_inst.ii3.i.ydata[25] ),
    .A2(_0439_),
    .B1(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0017_));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(net119),
    .B(\tokenflow_inst.i2.cg3.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0030_));
 sky130_fd_sc_hd__a21o_1 _0999_ (.A1(\tokenflow_inst.i10.d0.inv_chain[1] ),
    .A2(\tokenflow_inst.i10.cg.q ),
    .B1(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1000_ (.A(net127),
    .B(\tokenflow_inst.i8.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__a21o_1 _1001_ (.A1(net35),
    .A2(\tokenflow_inst.i8.ydata[53] ),
    .B1(\tokenflow_inst.i8.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__nand3_1 _1002_ (.A(net35),
    .B(\tokenflow_inst.i8.ydata[53] ),
    .C(\tokenflow_inst.i8.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0442_));
 sky130_fd_sc_hd__and3_1 _1003_ (.A(net127),
    .B(_0441_),
    .C(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__and3_1 _1004_ (.A(net35),
    .B(\tokenflow_inst.i8.ydata[54] ),
    .C(\tokenflow_inst.i8.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__a21oi_1 _1005_ (.A1(net35),
    .A2(\tokenflow_inst.i8.ydata[54] ),
    .B1(\tokenflow_inst.i8.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0444_));
 sky130_fd_sc_hd__o21ai_1 _1006_ (.A1(_0443_),
    .A2(_0444_),
    .B1(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0445_));
 sky130_fd_sc_hd__o311a_1 _1007_ (.A1(_0442_),
    .A2(_0443_),
    .A3(_0444_),
    .B1(_0445_),
    .C1(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__o21ba_1 _1008_ (.A1(_0442_),
    .A2(_0444_),
    .B1_N(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__a21oi_1 _1009_ (.A1(net35),
    .A2(\tokenflow_inst.i8.ydata[55] ),
    .B1(\tokenflow_inst.i8.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0447_));
 sky130_fd_sc_hd__and3_1 _1010_ (.A(net36),
    .B(\tokenflow_inst.i8.ydata[55] ),
    .C(\tokenflow_inst.i8.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__or2_1 _1011_ (.A(_0447_),
    .B(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__nand2_1 _1012_ (.A(_0446_),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_1 _1013_ (.A(_0446_),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__and3_1 _1014_ (.A(net125),
    .B(_0450_),
    .C(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__a21oi_1 _1015_ (.A1(net35),
    .A2(\tokenflow_inst.i8.ydata[56] ),
    .B1(\tokenflow_inst.i8.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0452_));
 sky130_fd_sc_hd__and3_1 _1016_ (.A(net35),
    .B(\tokenflow_inst.i8.ydata[56] ),
    .C(\tokenflow_inst.i8.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(_0452_),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0454_));
 sky130_fd_sc_hd__nand3b_1 _1018_ (.A_N(_0448_),
    .B(_0451_),
    .C(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0455_));
 sky130_fd_sc_hd__or3_2 _1019_ (.A(_0446_),
    .B(_0449_),
    .C(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0456_));
 sky130_fd_sc_hd__or3b_1 _1020_ (.A(_0452_),
    .B(_0453_),
    .C_N(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0457_));
 sky130_fd_sc_hd__and4_1 _1021_ (.A(net125),
    .B(_0455_),
    .C(_0456_),
    .D(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__and2b_1 _1022_ (.A_N(_0453_),
    .B(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__a21oi_1 _1023_ (.A1(net35),
    .A2(\tokenflow_inst.i8.ydata[57] ),
    .B1(\tokenflow_inst.i8.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0459_));
 sky130_fd_sc_hd__and3_1 _1024_ (.A(net35),
    .B(\tokenflow_inst.i8.ydata[57] ),
    .C(\tokenflow_inst.i8.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _1025_ (.A(_0459_),
    .B(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0461_));
 sky130_fd_sc_hd__a21oi_1 _1026_ (.A1(_0456_),
    .A2(_0458_),
    .B1(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0462_));
 sky130_fd_sc_hd__a31o_1 _1027_ (.A1(_0456_),
    .A2(_0458_),
    .A3(_0461_),
    .B1(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_1 _1028_ (.A(_0462_),
    .B(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0248_));
 sky130_fd_sc_hd__and3_1 _1029_ (.A(net34),
    .B(\tokenflow_inst.i8.ydata[58] ),
    .C(\tokenflow_inst.i8.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0464_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0465_));
 sky130_fd_sc_hd__a21oi_1 _1031_ (.A1(net34),
    .A2(\tokenflow_inst.i8.ydata[58] ),
    .B1(\tokenflow_inst.i8.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _1032_ (.A(_0464_),
    .B(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0467_));
 sky130_fd_sc_hd__or3_1 _1033_ (.A(_0460_),
    .B(_0462_),
    .C(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0468_));
 sky130_fd_sc_hd__o21ai_1 _1034_ (.A1(_0460_),
    .A2(_0462_),
    .B1(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0469_));
 sky130_fd_sc_hd__and3_1 _1035_ (.A(net114),
    .B(_0468_),
    .C(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__a21oi_1 _1036_ (.A1(net34),
    .A2(\tokenflow_inst.i8.ydata[59] ),
    .B1(\tokenflow_inst.i8.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0470_));
 sky130_fd_sc_hd__and3_1 _1037_ (.A(net34),
    .B(\tokenflow_inst.i8.ydata[7] ),
    .C(\tokenflow_inst.i8.ydata[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0471_));
 sky130_fd_sc_hd__or2_1 _1038_ (.A(_0470_),
    .B(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0472_));
 sky130_fd_sc_hd__and3_1 _1039_ (.A(_0465_),
    .B(_0469_),
    .C(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0473_));
 sky130_fd_sc_hd__a21oi_1 _1040_ (.A1(_0465_),
    .A2(_0469_),
    .B1(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0474_));
 sky130_fd_sc_hd__nor3_1 _1041_ (.A(net88),
    .B(_0473_),
    .C(_0474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0268_));
 sky130_fd_sc_hd__and3_1 _1042_ (.A(net34),
    .B(\tokenflow_inst.i8.ydata[60] ),
    .C(\tokenflow_inst.i8.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0475_));
 sky130_fd_sc_hd__a21oi_1 _1043_ (.A1(net34),
    .A2(\tokenflow_inst.i8.ydata[60] ),
    .B1(\tokenflow_inst.i8.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0476_));
 sky130_fd_sc_hd__a21o_1 _1044_ (.A1(net34),
    .A2(\tokenflow_inst.i8.ydata[60] ),
    .B1(\tokenflow_inst.i8.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _1045_ (.A(_0475_),
    .B(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0478_));
 sky130_fd_sc_hd__o21ai_1 _1046_ (.A1(_0471_),
    .A2(_0474_),
    .B1(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0479_));
 sky130_fd_sc_hd__or3_1 _1047_ (.A(_0471_),
    .B(_0474_),
    .C(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0480_));
 sky130_fd_sc_hd__and3_1 _1048_ (.A(net113),
    .B(_0479_),
    .C(_0480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__or4_1 _1049_ (.A(_0470_),
    .B(_0471_),
    .C(_0475_),
    .D(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0481_));
 sky130_fd_sc_hd__or3_1 _1050_ (.A(_0461_),
    .B(_0464_),
    .C(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0482_));
 sky130_fd_sc_hd__a211o_1 _1051_ (.A1(_0456_),
    .A2(_0458_),
    .B1(_0481_),
    .C1(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__and2b_1 _1052_ (.A_N(_0466_),
    .B(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0484_));
 sky130_fd_sc_hd__o21ba_1 _1053_ (.A1(_0464_),
    .A2(_0484_),
    .B1_N(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0485_));
 sky130_fd_sc_hd__a211oi_1 _1054_ (.A1(_0471_),
    .A2(_0477_),
    .B1(_0485_),
    .C1(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0486_));
 sky130_fd_sc_hd__and2_1 _1055_ (.A(_0483_),
    .B(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0487_));
 sky130_fd_sc_hd__a21oi_1 _1056_ (.A1(net33),
    .A2(\tokenflow_inst.i8.ydata[61] ),
    .B1(\tokenflow_inst.i8.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0488_));
 sky130_fd_sc_hd__and3_1 _1057_ (.A(\tokenflow_inst.i8.ydata[26] ),
    .B(\tokenflow_inst.i8.ydata[9] ),
    .C(\tokenflow_inst.i8.ydata[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0489_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0490_));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(_0488_),
    .B(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_1 _1060_ (.A(_0487_),
    .B(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0492_));
 sky130_fd_sc_hd__or2_1 _1061_ (.A(_0487_),
    .B(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0493_));
 sky130_fd_sc_hd__and3_1 _1062_ (.A(net99),
    .B(_0492_),
    .C(_0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _1063_ (.A(net31),
    .B(\tokenflow_inst.i8.ydata[62] ),
    .C(\tokenflow_inst.i8.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0494_));
 sky130_fd_sc_hd__a21oi_1 _1064_ (.A1(net31),
    .A2(\tokenflow_inst.i8.ydata[62] ),
    .B1(\tokenflow_inst.i8.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0495_));
 sky130_fd_sc_hd__or2_1 _1065_ (.A(_0494_),
    .B(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0496_));
 sky130_fd_sc_hd__nand3_1 _1066_ (.A(_0490_),
    .B(_0493_),
    .C(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0497_));
 sky130_fd_sc_hd__a21o_1 _1067_ (.A1(_0490_),
    .A2(_0493_),
    .B1(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0498_));
 sky130_fd_sc_hd__and3_1 _1068_ (.A(net99),
    .B(_0497_),
    .C(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__a21oi_1 _1069_ (.A1(net31),
    .A2(\tokenflow_inst.i8.ydata[63] ),
    .B1(\tokenflow_inst.i8.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0499_));
 sky130_fd_sc_hd__and3_1 _1070_ (.A(net31),
    .B(\tokenflow_inst.i8.ydata[11] ),
    .C(\tokenflow_inst.i8.ydata[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _1071_ (.A(_0499_),
    .B(_0500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0501_));
 sky130_fd_sc_hd__and2b_1 _1072_ (.A_N(_0494_),
    .B(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(_0501_),
    .B(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _1074_ (.A(_0501_),
    .B(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0504_));
 sky130_fd_sc_hd__and3b_1 _1075_ (.A_N(_0504_),
    .B(net94),
    .C(_0503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__and3_1 _1076_ (.A(net31),
    .B(\tokenflow_inst.i8.ydata[64] ),
    .C(\tokenflow_inst.i8.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _1077_ (.A1(net31),
    .A2(\tokenflow_inst.i8.ydata[64] ),
    .B1(\tokenflow_inst.i8.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0506_));
 sky130_fd_sc_hd__a21o_1 _1078_ (.A1(net31),
    .A2(\tokenflow_inst.i8.ydata[64] ),
    .B1(\tokenflow_inst.i8.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_1 _1079_ (.A(_0505_),
    .B(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0508_));
 sky130_fd_sc_hd__o21ai_1 _1080_ (.A1(_0500_),
    .A2(_0504_),
    .B1(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0509_));
 sky130_fd_sc_hd__or3_1 _1081_ (.A(_0500_),
    .B(_0504_),
    .C(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0510_));
 sky130_fd_sc_hd__and3_1 _1082_ (.A(net94),
    .B(_0509_),
    .C(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__a21oi_1 _1083_ (.A1(net32),
    .A2(\tokenflow_inst.i8.ydata[65] ),
    .B1(\tokenflow_inst.i8.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0511_));
 sky130_fd_sc_hd__and3_1 _1084_ (.A(net31),
    .B(\tokenflow_inst.i8.ydata[13] ),
    .C(\tokenflow_inst.i8.ydata[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _1085_ (.A(_0511_),
    .B(_0512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0513_));
 sky130_fd_sc_hd__or4_1 _1086_ (.A(_0499_),
    .B(_0500_),
    .C(_0505_),
    .D(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0514_));
 sky130_fd_sc_hd__or3_1 _1087_ (.A(_0491_),
    .B(_0496_),
    .C(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0515_));
 sky130_fd_sc_hd__and2b_1 _1088_ (.A_N(_0495_),
    .B(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0516_));
 sky130_fd_sc_hd__o21ba_1 _1089_ (.A1(_0494_),
    .A2(_0516_),
    .B1_N(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0517_));
 sky130_fd_sc_hd__a211oi_1 _1090_ (.A1(_0500_),
    .A2(_0507_),
    .B1(_0517_),
    .C1(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0518_));
 sky130_fd_sc_hd__o21a_1 _1091_ (.A1(_0487_),
    .A2(_0515_),
    .B1(_0518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0519_));
 sky130_fd_sc_hd__nand2_1 _1092_ (.A(_0513_),
    .B(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0520_));
 sky130_fd_sc_hd__or2_1 _1093_ (.A(_0513_),
    .B(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0522_));
 sky130_fd_sc_hd__and3_1 _1095_ (.A(net108),
    .B(_0520_),
    .C(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__a21oi_1 _1096_ (.A1(net31),
    .A2(\tokenflow_inst.i8.ydata[66] ),
    .B1(\tokenflow_inst.i8.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0523_));
 sky130_fd_sc_hd__and3_1 _1097_ (.A(net31),
    .B(\tokenflow_inst.i8.ydata[66] ),
    .C(\tokenflow_inst.i8.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0524_));
 sky130_fd_sc_hd__nor2_1 _1098_ (.A(_0523_),
    .B(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0525_));
 sky130_fd_sc_hd__and2b_1 _1099_ (.A_N(_0521_),
    .B(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0526_));
 sky130_fd_sc_hd__or3_1 _1100_ (.A(_0512_),
    .B(_0522_),
    .C(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_1 _1101_ (.A(_0512_),
    .B(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0528_));
 sky130_fd_sc_hd__and4b_1 _1102_ (.A_N(_0526_),
    .B(_0527_),
    .C(_0528_),
    .D(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__and3_1 _1103_ (.A(net33),
    .B(\tokenflow_inst.i8.ydata[15] ),
    .C(\tokenflow_inst.i8.ydata[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _1104_ (.A1(net33),
    .A2(\tokenflow_inst.i8.ydata[67] ),
    .B1(\tokenflow_inst.i8.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _1105_ (.A(_0529_),
    .B(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0531_));
 sky130_fd_sc_hd__a21o_1 _1106_ (.A1(_0512_),
    .A2(_0525_),
    .B1(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0532_));
 sky130_fd_sc_hd__o21a_1 _1107_ (.A1(_0526_),
    .A2(_0532_),
    .B1(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0533_));
 sky130_fd_sc_hd__nor2_1 _1108_ (.A(net89),
    .B(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0534_));
 sky130_fd_sc_hd__o31a_1 _1109_ (.A1(_0526_),
    .A2(_0531_),
    .A3(_0532_),
    .B1(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__a21oi_1 _1110_ (.A1(net33),
    .A2(\tokenflow_inst.i8.ydata[68] ),
    .B1(\tokenflow_inst.i8.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0535_));
 sky130_fd_sc_hd__and3_1 _1111_ (.A(net33),
    .B(\tokenflow_inst.i8.ydata[68] ),
    .C(\tokenflow_inst.i8.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(_0535_),
    .B(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0537_));
 sky130_fd_sc_hd__or3_1 _1113_ (.A(_0529_),
    .B(_0533_),
    .C(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0538_));
 sky130_fd_sc_hd__o21ai_1 _1114_ (.A1(_0529_),
    .A2(_0533_),
    .B1(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0539_));
 sky130_fd_sc_hd__and3_1 _1115_ (.A(net108),
    .B(_0538_),
    .C(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__and4b_1 _1116_ (.A_N(_0513_),
    .B(_0525_),
    .C(_0531_),
    .D(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _1117_ (.A(_0540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _1118_ (.A(_0529_),
    .B(_0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0542_));
 sky130_fd_sc_hd__or3_1 _1119_ (.A(_0530_),
    .B(_0535_),
    .C(_0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0543_));
 sky130_fd_sc_hd__o21ba_1 _1120_ (.A1(_0518_),
    .A2(_0541_),
    .B1_N(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0544_));
 sky130_fd_sc_hd__a211o_1 _1121_ (.A1(_0483_),
    .A2(_0486_),
    .B1(_0515_),
    .C1(_0541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0545_));
 sky130_fd_sc_hd__and3_1 _1122_ (.A(_0543_),
    .B(_0544_),
    .C(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0546_));
 sky130_fd_sc_hd__a21o_1 _1123_ (.A1(net36),
    .A2(\tokenflow_inst.i8.ydata[69] ),
    .B1(\tokenflow_inst.i8.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0547_));
 sky130_fd_sc_hd__nand3_1 _1124_ (.A(net34),
    .B(\tokenflow_inst.i8.ydata[17] ),
    .C(\tokenflow_inst.i8.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _1125_ (.A(_0547_),
    .B(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(_0546_),
    .B(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0550_));
 sky130_fd_sc_hd__a31o_1 _1127_ (.A1(_0543_),
    .A2(_0544_),
    .A3(_0545_),
    .B1(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _1128_ (.A(net108),
    .B(_0550_),
    .C(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _1129_ (.A1(net36),
    .A2(\tokenflow_inst.i8.ydata[70] ),
    .B1(\tokenflow_inst.i8.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0552_));
 sky130_fd_sc_hd__and3_1 _1130_ (.A(net36),
    .B(\tokenflow_inst.i8.ydata[18] ),
    .C(\tokenflow_inst.i8.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _1131_ (.A(_0552_),
    .B(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0554_));
 sky130_fd_sc_hd__and3_1 _1132_ (.A(_0548_),
    .B(_0551_),
    .C(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(_0551_),
    .B(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(_0548_),
    .B(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0557_));
 sky130_fd_sc_hd__nor4_1 _1135_ (.A(net88),
    .B(_0555_),
    .C(_0556_),
    .D(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0206_));
 sky130_fd_sc_hd__a21o_1 _1136_ (.A1(net36),
    .A2(\tokenflow_inst.i8.ydata[71] ),
    .B1(\tokenflow_inst.i8.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0558_));
 sky130_fd_sc_hd__nand3_1 _1137_ (.A(net35),
    .B(\tokenflow_inst.i8.ydata[19] ),
    .C(\tokenflow_inst.i8.ydata[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(_0558_),
    .B(_0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0560_));
 sky130_fd_sc_hd__nor2_1 _1139_ (.A(_0553_),
    .B(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(_0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0562_));
 sky130_fd_sc_hd__or3b_1 _1141_ (.A(_0556_),
    .B(_0562_),
    .C_N(_0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0563_));
 sky130_fd_sc_hd__o21bai_1 _1142_ (.A1(_0556_),
    .A2(_0562_),
    .B1_N(_0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0564_));
 sky130_fd_sc_hd__and3_1 _1143_ (.A(net123),
    .B(_0563_),
    .C(_0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _1144_ (.A(net34),
    .B(\tokenflow_inst.i8.ydata[72] ),
    .C(\tokenflow_inst.i8.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0565_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(_0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1146_ (.A1(net34),
    .A2(\tokenflow_inst.i8.ydata[72] ),
    .B1(\tokenflow_inst.i8.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0567_));
 sky130_fd_sc_hd__or2_1 _1147_ (.A(_0565_),
    .B(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_1 _1148_ (.A1(_0559_),
    .A2(_0564_),
    .B1(_0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _1149_ (.A(net123),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0570_));
 sky130_fd_sc_hd__a31oi_1 _1150_ (.A1(_0559_),
    .A2(_0564_),
    .A3(_0568_),
    .B1(_0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0209_));
 sky130_fd_sc_hd__or2_1 _1151_ (.A(_0560_),
    .B(_0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0571_));
 sky130_fd_sc_hd__o221a_1 _1152_ (.A1(_0559_),
    .A2(_0567_),
    .B1(_0571_),
    .B2(_0561_),
    .C1(_0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0572_));
 sky130_fd_sc_hd__o31a_2 _1153_ (.A1(_0551_),
    .A2(_0554_),
    .A3(_0571_),
    .B1(_0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0573_));
 sky130_fd_sc_hd__a21o_1 _1154_ (.A1(net33),
    .A2(\tokenflow_inst.i8.ydata[73] ),
    .B1(\tokenflow_inst.i8.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0574_));
 sky130_fd_sc_hd__nand3_1 _1155_ (.A(net33),
    .B(\tokenflow_inst.i8.ydata[21] ),
    .C(\tokenflow_inst.i8.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1156_ (.A(_0574_),
    .B(_0575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0576_));
 sky130_fd_sc_hd__o21ai_1 _1157_ (.A1(_0573_),
    .A2(_0576_),
    .B1(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0577_));
 sky130_fd_sc_hd__a21oi_1 _1158_ (.A1(_0573_),
    .A2(_0576_),
    .B1(_0577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0210_));
 sky130_fd_sc_hd__a21oi_1 _1159_ (.A1(net33),
    .A2(\tokenflow_inst.i8.ydata[74] ),
    .B1(\tokenflow_inst.i8.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0578_));
 sky130_fd_sc_hd__and3_1 _1160_ (.A(net33),
    .B(\tokenflow_inst.i8.ydata[22] ),
    .C(\tokenflow_inst.i8.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0579_));
 sky130_fd_sc_hd__or2_1 _1161_ (.A(_0578_),
    .B(_0579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0580_));
 sky130_fd_sc_hd__o211ai_1 _1162_ (.A1(_0573_),
    .A2(_0576_),
    .B1(_0580_),
    .C1(_0575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0581_));
 sky130_fd_sc_hd__or3_1 _1163_ (.A(_0573_),
    .B(_0576_),
    .C(_0580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0582_));
 sky130_fd_sc_hd__o2111a_1 _1164_ (.A1(_0575_),
    .A2(_0580_),
    .B1(_0581_),
    .C1(_0582_),
    .D1(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__o21ba_1 _1165_ (.A1(_0575_),
    .A2(_0578_),
    .B1_N(_0579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0583_));
 sky130_fd_sc_hd__o31ai_2 _1166_ (.A1(_0573_),
    .A2(_0576_),
    .A3(_0580_),
    .B1(_0583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0584_));
 sky130_fd_sc_hd__a21oi_1 _1167_ (.A1(net32),
    .A2(\tokenflow_inst.i8.ydata[75] ),
    .B1(\tokenflow_inst.i8.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0585_));
 sky130_fd_sc_hd__and3_1 _1168_ (.A(net32),
    .B(\tokenflow_inst.i8.ydata[23] ),
    .C(\tokenflow_inst.i8.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0586_));
 sky130_fd_sc_hd__nor2_1 _1169_ (.A(_0585_),
    .B(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0587_));
 sky130_fd_sc_hd__a21oi_1 _1170_ (.A1(_0584_),
    .A2(_0587_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0588_));
 sky130_fd_sc_hd__o21a_1 _1171_ (.A1(_0584_),
    .A2(_0587_),
    .B1(_0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__a21oi_1 _1172_ (.A1(net32),
    .A2(\tokenflow_inst.i8.ydata[76] ),
    .B1(\tokenflow_inst.i8.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0589_));
 sky130_fd_sc_hd__and3_1 _1173_ (.A(net32),
    .B(\tokenflow_inst.i8.ydata[24] ),
    .C(\tokenflow_inst.i8.ydata[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0590_));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _1175_ (.A(_0589_),
    .B(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0592_));
 sky130_fd_sc_hd__a211o_1 _1176_ (.A1(_0584_),
    .A2(_0587_),
    .B1(_0592_),
    .C1(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0593_));
 sky130_fd_sc_hd__nand3_1 _1177_ (.A(_0584_),
    .B(_0587_),
    .C(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0586_),
    .B(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0595_));
 sky130_fd_sc_hd__and4_1 _1179_ (.A(net104),
    .B(_0593_),
    .C(_0594_),
    .D(_0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(net32),
    .B(\tokenflow_inst.i8.ydata[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0596_));
 sky130_fd_sc_hd__xor2_1 _1181_ (.A(\tokenflow_inst.i8.ydata[25] ),
    .B(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0597_));
 sky130_fd_sc_hd__a31o_1 _1182_ (.A1(_0591_),
    .A2(_0594_),
    .A3(_0595_),
    .B1(_0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0598_));
 sky130_fd_sc_hd__a41o_1 _1183_ (.A1(_0591_),
    .A2(_0594_),
    .A3(_0595_),
    .A4(_0597_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0599_));
 sky130_fd_sc_hd__and2b_1 _1184_ (.A_N(_0599_),
    .B(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__and2_1 _1185_ (.A(net116),
    .B(\tokenflow_inst.i8.ydata[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _1186_ (.A(net145),
    .B(\tokenflow_inst.i8.ydata[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _1187_ (.A(net116),
    .B(\tokenflow_inst.i8.ydata[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__and2_1 _1188_ (.A(net116),
    .B(\tokenflow_inst.i8.ydata[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__and2_1 _1189_ (.A(net145),
    .B(\tokenflow_inst.i8.ydata[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__and2_1 _1190_ (.A(net112),
    .B(\tokenflow_inst.i8.ydata[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(net111),
    .B(\tokenflow_inst.i8.ydata[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__and2_1 _1192_ (.A(net110),
    .B(\tokenflow_inst.i8.ydata[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__and2_1 _1193_ (.A(net112),
    .B(\tokenflow_inst.i8.ydata[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__and2_1 _1194_ (.A(net97),
    .B(\tokenflow_inst.i8.ydata[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__and2_1 _1195_ (.A(net91),
    .B(\tokenflow_inst.i8.ydata[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__and2_1 _1196_ (.A(net91),
    .B(\tokenflow_inst.i8.ydata[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__and2_1 _1197_ (.A(net90),
    .B(\tokenflow_inst.i8.ydata[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _1198_ (.A(net90),
    .B(\tokenflow_inst.i8.ydata[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__and2_1 _1199_ (.A(net92),
    .B(\tokenflow_inst.i8.ydata[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__and2_1 _1200_ (.A(net92),
    .B(\tokenflow_inst.i8.ydata[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(net96),
    .B(\tokenflow_inst.i8.ydata[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__and2_1 _1202_ (.A(net97),
    .B(\tokenflow_inst.i8.ydata[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _1203_ (.A(net110),
    .B(\tokenflow_inst.i8.ydata[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _1204_ (.A(net110),
    .B(\tokenflow_inst.i8.ydata[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _1205_ (.A(net98),
    .B(\tokenflow_inst.i8.ydata[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__and2_1 _1206_ (.A(net97),
    .B(\tokenflow_inst.i8.ydata[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__and2_1 _1207_ (.A(net96),
    .B(\tokenflow_inst.i8.ydata[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _1208_ (.A(net93),
    .B(\tokenflow_inst.i8.ydata[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__and2_1 _1209_ (.A(net127),
    .B(\tokenflow_inst.i8.ydata[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _1210_ (.A(net127),
    .B(\tokenflow_inst.i8.ydata[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__and2_1 _1211_ (.A(net125),
    .B(\tokenflow_inst.i8.ydata[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _1212_ (.A(net125),
    .B(\tokenflow_inst.i8.ydata[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__and2_1 _1213_ (.A(net117),
    .B(\tokenflow_inst.i8.ydata[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__and2_1 _1214_ (.A(net114),
    .B(\tokenflow_inst.i8.ydata[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__and2_1 _1215_ (.A(net113),
    .B(\tokenflow_inst.i8.ydata[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__and2_1 _1216_ (.A(net113),
    .B(\tokenflow_inst.i8.ydata[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(net99),
    .B(\tokenflow_inst.i8.ydata[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _1218_ (.A(net101),
    .B(\tokenflow_inst.i8.ydata[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__and2_1 _1219_ (.A(net95),
    .B(\tokenflow_inst.i8.ydata[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__and2_1 _1220_ (.A(net102),
    .B(\tokenflow_inst.i8.ydata[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__and2_1 _1221_ (.A(net102),
    .B(\tokenflow_inst.i8.ydata[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__and2_1 _1222_ (.A(net102),
    .B(\tokenflow_inst.i8.ydata[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(net108),
    .B(\tokenflow_inst.i8.ydata[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _1224_ (.A(net106),
    .B(\tokenflow_inst.i8.ydata[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__and2_1 _1225_ (.A(net122),
    .B(\tokenflow_inst.i8.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__and2_1 _1226_ (.A(net123),
    .B(\tokenflow_inst.i8.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__and2_1 _1227_ (.A(net123),
    .B(\tokenflow_inst.i8.ydata[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__and2_1 _1228_ (.A(net123),
    .B(\tokenflow_inst.i8.ydata[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(net106),
    .B(\tokenflow_inst.i8.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _1230_ (.A(net106),
    .B(\tokenflow_inst.i8.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _1231_ (.A(net104),
    .B(\tokenflow_inst.i8.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__and2_1 _1232_ (.A(net104),
    .B(\tokenflow_inst.i8.ydata[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__a21o_1 _1233_ (.A1(net63),
    .A2(\tokenflow_inst.i6.ydata[52] ),
    .B1(\tokenflow_inst.i6.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0600_));
 sky130_fd_sc_hd__nand3_1 _1234_ (.A(net63),
    .B(\tokenflow_inst.i6.ydata[52] ),
    .C(\tokenflow_inst.i6.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0601_));
 sky130_fd_sc_hd__and3_1 _1235_ (.A(net127),
    .B(_0600_),
    .C(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__and3_1 _1236_ (.A(net63),
    .B(\tokenflow_inst.i6.ydata[53] ),
    .C(\tokenflow_inst.i6.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0602_));
 sky130_fd_sc_hd__a21oi_1 _1237_ (.A1(net63),
    .A2(\tokenflow_inst.i6.ydata[53] ),
    .B1(\tokenflow_inst.i6.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0603_));
 sky130_fd_sc_hd__o21ai_1 _1238_ (.A1(_0602_),
    .A2(_0603_),
    .B1(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0604_));
 sky130_fd_sc_hd__o311a_1 _1239_ (.A1(_0601_),
    .A2(_0602_),
    .A3(_0603_),
    .B1(_0604_),
    .C1(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__o21ba_1 _1240_ (.A1(_0601_),
    .A2(_0603_),
    .B1_N(_0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0605_));
 sky130_fd_sc_hd__a21oi_1 _1241_ (.A1(net63),
    .A2(\tokenflow_inst.i6.ydata[54] ),
    .B1(\tokenflow_inst.i6.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0606_));
 sky130_fd_sc_hd__and3_1 _1242_ (.A(net63),
    .B(\tokenflow_inst.i6.ydata[54] ),
    .C(\tokenflow_inst.i6.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0607_));
 sky130_fd_sc_hd__or2_1 _1243_ (.A(_0606_),
    .B(_0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _1244_ (.A(_0605_),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0609_));
 sky130_fd_sc_hd__a21o_1 _1245_ (.A1(_0605_),
    .A2(_0608_),
    .B1(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_1 _1246_ (.A(_0609_),
    .B(_0610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0296_));
 sky130_fd_sc_hd__a21o_1 _1247_ (.A1(net63),
    .A2(\tokenflow_inst.i6.ydata[55] ),
    .B1(\tokenflow_inst.i6.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0611_));
 sky130_fd_sc_hd__nand3_1 _1248_ (.A(net63),
    .B(\tokenflow_inst.i6.ydata[55] ),
    .C(\tokenflow_inst.i6.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0612_));
 sky130_fd_sc_hd__and2_1 _1249_ (.A(_0611_),
    .B(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0613_));
 sky130_fd_sc_hd__or3b_2 _1250_ (.A(_0605_),
    .B(_0608_),
    .C_N(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0614_));
 sky130_fd_sc_hd__or3_1 _1251_ (.A(_0607_),
    .B(_0609_),
    .C(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0607_),
    .B(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0616_));
 sky130_fd_sc_hd__and4_1 _1253_ (.A(net125),
    .B(_0614_),
    .C(_0615_),
    .D(_0616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__a21boi_1 _1254_ (.A1(_0607_),
    .A2(_0611_),
    .B1_N(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0617_));
 sky130_fd_sc_hd__a21oi_1 _1255_ (.A1(net63),
    .A2(\tokenflow_inst.i6.ydata[56] ),
    .B1(\tokenflow_inst.i6.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0618_));
 sky130_fd_sc_hd__and3_1 _1256_ (.A(net63),
    .B(\tokenflow_inst.i6.ydata[56] ),
    .C(\tokenflow_inst.i6.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _1257_ (.A(_0618_),
    .B(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0620_));
 sky130_fd_sc_hd__a21oi_1 _1258_ (.A1(_0614_),
    .A2(_0617_),
    .B1(_0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0621_));
 sky130_fd_sc_hd__a31o_1 _1259_ (.A1(_0614_),
    .A2(_0617_),
    .A3(_0620_),
    .B1(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _1260_ (.A(_0621_),
    .B(_0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0318_));
 sky130_fd_sc_hd__and3_1 _1261_ (.A(net61),
    .B(\tokenflow_inst.i6.ydata[57] ),
    .C(\tokenflow_inst.i6.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0623_));
 sky130_fd_sc_hd__inv_2 _1262_ (.A(_0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0624_));
 sky130_fd_sc_hd__a21oi_1 _1263_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[57] ),
    .B1(\tokenflow_inst.i6.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0625_));
 sky130_fd_sc_hd__nor2_1 _1264_ (.A(_0623_),
    .B(_0625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0626_));
 sky130_fd_sc_hd__or3_1 _1265_ (.A(_0619_),
    .B(_0621_),
    .C(_0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0627_));
 sky130_fd_sc_hd__o21ai_1 _1266_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0628_));
 sky130_fd_sc_hd__and3_1 _1267_ (.A(net122),
    .B(_0627_),
    .C(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__a21oi_1 _1268_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[58] ),
    .B1(\tokenflow_inst.i6.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0629_));
 sky130_fd_sc_hd__and3_1 _1269_ (.A(net61),
    .B(\tokenflow_inst.i6.ydata[6] ),
    .C(\tokenflow_inst.i6.ydata[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0630_));
 sky130_fd_sc_hd__or2_1 _1270_ (.A(_0629_),
    .B(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _1271_ (.A(_0624_),
    .B(_0628_),
    .C(_0631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0632_));
 sky130_fd_sc_hd__a21oi_1 _1272_ (.A1(_0624_),
    .A2(_0628_),
    .B1(_0631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0633_));
 sky130_fd_sc_hd__nor3_1 _1273_ (.A(net88),
    .B(_0632_),
    .C(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0338_));
 sky130_fd_sc_hd__and3_1 _1274_ (.A(net61),
    .B(\tokenflow_inst.i6.ydata[59] ),
    .C(\tokenflow_inst.i6.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0634_));
 sky130_fd_sc_hd__a21oi_1 _1275_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[59] ),
    .B1(\tokenflow_inst.i6.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0635_));
 sky130_fd_sc_hd__a21o_1 _1276_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[59] ),
    .B1(\tokenflow_inst.i6.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0636_));
 sky130_fd_sc_hd__nor2_1 _1277_ (.A(_0634_),
    .B(_0635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0637_));
 sky130_fd_sc_hd__o21ai_1 _1278_ (.A1(_0630_),
    .A2(_0633_),
    .B1(_0637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0638_));
 sky130_fd_sc_hd__or3_1 _1279_ (.A(_0630_),
    .B(_0633_),
    .C(_0637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _1280_ (.A(net122),
    .B(_0638_),
    .C(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__or4_1 _1281_ (.A(_0629_),
    .B(_0630_),
    .C(_0634_),
    .D(_0635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0640_));
 sky130_fd_sc_hd__or3_1 _1282_ (.A(_0620_),
    .B(_0623_),
    .C(_0625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0641_));
 sky130_fd_sc_hd__a211o_1 _1283_ (.A1(_0614_),
    .A2(_0617_),
    .B1(_0640_),
    .C1(_0641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0642_));
 sky130_fd_sc_hd__and2b_1 _1284_ (.A_N(_0625_),
    .B(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0643_));
 sky130_fd_sc_hd__o21ba_1 _1285_ (.A1(_0623_),
    .A2(_0643_),
    .B1_N(_0640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0644_));
 sky130_fd_sc_hd__a211oi_1 _1286_ (.A1(_0630_),
    .A2(_0636_),
    .B1(_0644_),
    .C1(_0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0645_));
 sky130_fd_sc_hd__and2_1 _1287_ (.A(_0642_),
    .B(_0645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0646_));
 sky130_fd_sc_hd__a21oi_1 _1288_ (.A1(net60),
    .A2(\tokenflow_inst.i6.ydata[60] ),
    .B1(\tokenflow_inst.i6.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0647_));
 sky130_fd_sc_hd__and3_1 _1289_ (.A(net60),
    .B(\tokenflow_inst.i6.ydata[8] ),
    .C(\tokenflow_inst.i6.ydata[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0648_));
 sky130_fd_sc_hd__or2_1 _1290_ (.A(_0647_),
    .B(_0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0649_));
 sky130_fd_sc_hd__nor2_1 _1291_ (.A(_0646_),
    .B(_0649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0650_));
 sky130_fd_sc_hd__a31o_1 _1292_ (.A1(_0642_),
    .A2(_0645_),
    .A3(_0649_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _1293_ (.A(_0650_),
    .B(_0651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0348_));
 sky130_fd_sc_hd__and3_1 _1294_ (.A(net60),
    .B(\tokenflow_inst.i6.ydata[61] ),
    .C(\tokenflow_inst.i6.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0652_));
 sky130_fd_sc_hd__inv_2 _1295_ (.A(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0653_));
 sky130_fd_sc_hd__a21oi_1 _1296_ (.A1(net60),
    .A2(\tokenflow_inst.i6.ydata[61] ),
    .B1(\tokenflow_inst.i6.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _1297_ (.A(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0655_));
 sky130_fd_sc_hd__or2_1 _1298_ (.A(_0652_),
    .B(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0656_));
 sky130_fd_sc_hd__or3b_1 _1299_ (.A(_0648_),
    .B(_0650_),
    .C_N(_0656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0657_));
 sky130_fd_sc_hd__o21bai_1 _1300_ (.A1(_0648_),
    .A2(_0650_),
    .B1_N(_0656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0658_));
 sky130_fd_sc_hd__and3_1 _1301_ (.A(net108),
    .B(_0657_),
    .C(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__a21oi_1 _1302_ (.A1(net59),
    .A2(\tokenflow_inst.i6.ydata[62] ),
    .B1(\tokenflow_inst.i6.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0659_));
 sky130_fd_sc_hd__and3_1 _1303_ (.A(net59),
    .B(\tokenflow_inst.i6.ydata[10] ),
    .C(\tokenflow_inst.i6.ydata[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0660_));
 sky130_fd_sc_hd__or2_1 _1304_ (.A(_0659_),
    .B(_0660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0661_));
 sky130_fd_sc_hd__and3_1 _1305_ (.A(_0653_),
    .B(_0658_),
    .C(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0662_));
 sky130_fd_sc_hd__a21oi_1 _1306_ (.A1(_0653_),
    .A2(_0658_),
    .B1(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0663_));
 sky130_fd_sc_hd__nor3_1 _1307_ (.A(net89),
    .B(_0662_),
    .C(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0275_));
 sky130_fd_sc_hd__and3_1 _1308_ (.A(net60),
    .B(\tokenflow_inst.i6.ydata[63] ),
    .C(\tokenflow_inst.i6.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0664_));
 sky130_fd_sc_hd__a21oi_1 _1309_ (.A1(net60),
    .A2(\tokenflow_inst.i6.ydata[63] ),
    .B1(\tokenflow_inst.i6.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0665_));
 sky130_fd_sc_hd__a21o_1 _1310_ (.A1(net60),
    .A2(\tokenflow_inst.i6.ydata[63] ),
    .B1(\tokenflow_inst.i6.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0666_));
 sky130_fd_sc_hd__nor2_1 _1311_ (.A(_0664_),
    .B(_0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0667_));
 sky130_fd_sc_hd__o21ai_1 _1312_ (.A1(_0660_),
    .A2(_0663_),
    .B1(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0668_));
 sky130_fd_sc_hd__or3_1 _1313_ (.A(_0660_),
    .B(_0663_),
    .C(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0669_));
 sky130_fd_sc_hd__and3_1 _1314_ (.A(net108),
    .B(_0668_),
    .C(_0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__a21oi_1 _1315_ (.A1(net59),
    .A2(\tokenflow_inst.i6.ydata[64] ),
    .B1(\tokenflow_inst.i6.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0670_));
 sky130_fd_sc_hd__and3_1 _1316_ (.A(net59),
    .B(\tokenflow_inst.i6.ydata[12] ),
    .C(\tokenflow_inst.i6.ydata[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0671_));
 sky130_fd_sc_hd__or2_1 _1317_ (.A(_0670_),
    .B(_0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0672_));
 sky130_fd_sc_hd__or3_1 _1318_ (.A(_0661_),
    .B(_0664_),
    .C(_0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0673_));
 sky130_fd_sc_hd__a21oi_1 _1319_ (.A1(_0648_),
    .A2(_0655_),
    .B1(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0674_));
 sky130_fd_sc_hd__a21oi_1 _1320_ (.A1(_0660_),
    .A2(_0666_),
    .B1(_0664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0675_));
 sky130_fd_sc_hd__o21a_1 _1321_ (.A1(_0673_),
    .A2(_0674_),
    .B1(_0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0676_));
 sky130_fd_sc_hd__or3_1 _1322_ (.A(_0649_),
    .B(_0656_),
    .C(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0677_));
 sky130_fd_sc_hd__o21a_1 _1323_ (.A1(_0646_),
    .A2(_0677_),
    .B1(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0678_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(_0672_),
    .B(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0679_));
 sky130_fd_sc_hd__or2_1 _1325_ (.A(_0672_),
    .B(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0680_));
 sky130_fd_sc_hd__and3_1 _1326_ (.A(net103),
    .B(_0679_),
    .C(_0680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _1327_ (.A1(net59),
    .A2(\tokenflow_inst.i6.ydata[65] ),
    .B1(\tokenflow_inst.i6.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0681_));
 sky130_fd_sc_hd__and3_1 _1328_ (.A(net59),
    .B(\tokenflow_inst.i6.ydata[65] ),
    .C(\tokenflow_inst.i6.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _1329_ (.A(_0681_),
    .B(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0683_));
 sky130_fd_sc_hd__or2_1 _1330_ (.A(_0681_),
    .B(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0684_));
 sky130_fd_sc_hd__nand3b_1 _1331_ (.A_N(_0671_),
    .B(_0680_),
    .C(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0685_));
 sky130_fd_sc_hd__or2_1 _1332_ (.A(_0680_),
    .B(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(_0671_),
    .B(_0683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0687_));
 sky130_fd_sc_hd__and4_1 _1334_ (.A(net103),
    .B(_0685_),
    .C(_0686_),
    .D(_0687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _1335_ (.A1(net58),
    .A2(\tokenflow_inst.i6.ydata[66] ),
    .B1(\tokenflow_inst.i6.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0688_));
 sky130_fd_sc_hd__nand3_1 _1336_ (.A(net59),
    .B(\tokenflow_inst.i6.ydata[14] ),
    .C(\tokenflow_inst.i6.ydata[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1337_ (.A(_0688_),
    .B(_0689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0690_));
 sky130_fd_sc_hd__a21oi_1 _1338_ (.A1(_0671_),
    .A2(_0683_),
    .B1(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0691_));
 sky130_fd_sc_hd__nand3_1 _1339_ (.A(_0686_),
    .B(_0690_),
    .C(_0691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0692_));
 sky130_fd_sc_hd__a21o_1 _1340_ (.A1(_0686_),
    .A2(_0691_),
    .B1(_0690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _1341_ (.A(net103),
    .B(_0692_),
    .C(_0693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__and3_1 _1342_ (.A(net58),
    .B(\tokenflow_inst.i6.ydata[67] ),
    .C(\tokenflow_inst.i6.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0694_));
 sky130_fd_sc_hd__a21oi_1 _1343_ (.A1(net58),
    .A2(\tokenflow_inst.i6.ydata[67] ),
    .B1(\tokenflow_inst.i6.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0695_));
 sky130_fd_sc_hd__a211o_1 _1344_ (.A1(_0689_),
    .A2(_0693_),
    .B1(_0694_),
    .C1(_0695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0696_));
 sky130_fd_sc_hd__o211ai_1 _1345_ (.A1(_0694_),
    .A2(_0695_),
    .B1(_0689_),
    .C1(_0693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0697_));
 sky130_fd_sc_hd__and3_1 _1346_ (.A(net103),
    .B(_0696_),
    .C(_0697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _1347_ (.A(net61),
    .B(\tokenflow_inst.i6.ydata[16] ),
    .C(\tokenflow_inst.i6.ydata[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0698_));
 sky130_fd_sc_hd__a21oi_1 _1348_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[68] ),
    .B1(\tokenflow_inst.i6.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0699_));
 sky130_fd_sc_hd__or2_1 _1349_ (.A(_0698_),
    .B(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0700_));
 sky130_fd_sc_hd__or3_1 _1350_ (.A(_0690_),
    .B(_0694_),
    .C(_0695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0701_));
 sky130_fd_sc_hd__or3_1 _1351_ (.A(_0672_),
    .B(_0684_),
    .C(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0702_));
 sky130_fd_sc_hd__o21ba_1 _1352_ (.A1(_0689_),
    .A2(_0695_),
    .B1_N(_0694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0703_));
 sky130_fd_sc_hd__o221a_1 _1353_ (.A1(_0691_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0676_),
    .C1(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0704_));
 sky130_fd_sc_hd__a211o_1 _1354_ (.A1(_0642_),
    .A2(_0645_),
    .B1(_0677_),
    .C1(_0702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0705_));
 sky130_fd_sc_hd__and2_1 _1355_ (.A(_0704_),
    .B(_0705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0706_));
 sky130_fd_sc_hd__nand2_1 _1356_ (.A(_0700_),
    .B(_0706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0707_));
 sky130_fd_sc_hd__nor2_1 _1357_ (.A(_0700_),
    .B(_0706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0708_));
 sky130_fd_sc_hd__and3b_1 _1358_ (.A_N(_0708_),
    .B(net108),
    .C(_0707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1359_ (.A1(net62),
    .A2(\tokenflow_inst.i6.ydata[69] ),
    .B1(\tokenflow_inst.i6.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0709_));
 sky130_fd_sc_hd__and3_1 _1360_ (.A(net62),
    .B(\tokenflow_inst.i6.ydata[17] ),
    .C(\tokenflow_inst.i6.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0710_));
 sky130_fd_sc_hd__nand3_1 _1361_ (.A(net62),
    .B(\tokenflow_inst.i6.ydata[17] ),
    .C(\tokenflow_inst.i6.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0711_));
 sky130_fd_sc_hd__nor2_1 _1362_ (.A(_0709_),
    .B(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0712_));
 sky130_fd_sc_hd__or3_1 _1363_ (.A(_0698_),
    .B(_0708_),
    .C(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0713_));
 sky130_fd_sc_hd__o21ai_1 _1364_ (.A1(_0698_),
    .A2(_0708_),
    .B1(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0714_));
 sky130_fd_sc_hd__and3_1 _1365_ (.A(net122),
    .B(_0713_),
    .C(_0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__a21oi_1 _1366_ (.A1(net64),
    .A2(\tokenflow_inst.i6.ydata[70] ),
    .B1(\tokenflow_inst.i6.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0715_));
 sky130_fd_sc_hd__and3_1 _1367_ (.A(net64),
    .B(\tokenflow_inst.i6.ydata[18] ),
    .C(\tokenflow_inst.i6.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0716_));
 sky130_fd_sc_hd__or2_1 _1368_ (.A(_0715_),
    .B(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0717_));
 sky130_fd_sc_hd__a21o_1 _1369_ (.A1(_0698_),
    .A2(_0712_),
    .B1(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0718_));
 sky130_fd_sc_hd__nand3_1 _1370_ (.A(_0711_),
    .B(_0714_),
    .C(_0717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _1371_ (.A1(_0711_),
    .A2(_0714_),
    .B1(_0717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0720_));
 sky130_fd_sc_hd__and3b_1 _1372_ (.A_N(_0720_),
    .B(net123),
    .C(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__and3_1 _1373_ (.A(net64),
    .B(\tokenflow_inst.i6.ydata[71] ),
    .C(\tokenflow_inst.i6.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _1374_ (.A1(net64),
    .A2(\tokenflow_inst.i6.ydata[71] ),
    .B1(\tokenflow_inst.i6.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0722_));
 sky130_fd_sc_hd__and2b_1 _1375_ (.A_N(_0721_),
    .B(_0722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0723_));
 sky130_fd_sc_hd__or3_1 _1376_ (.A(_0716_),
    .B(_0720_),
    .C(_0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0724_));
 sky130_fd_sc_hd__o21ai_1 _1377_ (.A1(_0716_),
    .A2(_0720_),
    .B1(_0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0725_));
 sky130_fd_sc_hd__and3_1 _1378_ (.A(net123),
    .B(_0724_),
    .C(_0725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__and2b_1 _1379_ (.A_N(_0717_),
    .B(_0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0726_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(_0712_),
    .B(_0726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0727_));
 sky130_fd_sc_hd__a211oi_2 _1381_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0727_),
    .C1(_0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0728_));
 sky130_fd_sc_hd__and2_1 _1382_ (.A(_0718_),
    .B(_0726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0729_));
 sky130_fd_sc_hd__a21o_1 _1383_ (.A1(_0716_),
    .A2(_0722_),
    .B1(_0721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0730_));
 sky130_fd_sc_hd__or3_1 _1384_ (.A(_0728_),
    .B(_0729_),
    .C(_0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0731_));
 sky130_fd_sc_hd__a21oi_1 _1385_ (.A1(net62),
    .A2(\tokenflow_inst.i6.ydata[72] ),
    .B1(\tokenflow_inst.i6.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0732_));
 sky130_fd_sc_hd__and3_1 _1386_ (.A(net62),
    .B(\tokenflow_inst.i6.ydata[20] ),
    .C(\tokenflow_inst.i6.ydata[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_2 _1387_ (.A(_0732_),
    .B(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _1388_ (.A1(_0731_),
    .A2(_0734_),
    .B1(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0735_));
 sky130_fd_sc_hd__o21a_1 _1389_ (.A1(_0731_),
    .A2(_0734_),
    .B1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__a21oi_1 _1390_ (.A1(net61),
    .A2(\tokenflow_inst.i6.ydata[73] ),
    .B1(\tokenflow_inst.i6.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0736_));
 sky130_fd_sc_hd__and3_1 _1391_ (.A(net62),
    .B(\tokenflow_inst.i6.ydata[21] ),
    .C(\tokenflow_inst.i6.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0737_));
 sky130_fd_sc_hd__nor2_2 _1392_ (.A(_0736_),
    .B(_0737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0738_));
 sky130_fd_sc_hd__a211o_1 _1393_ (.A1(_0731_),
    .A2(_0734_),
    .B1(_0738_),
    .C1(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0739_));
 sky130_fd_sc_hd__o311ai_4 _1394_ (.A1(_0728_),
    .A2(_0729_),
    .A3(_0730_),
    .B1(_0734_),
    .C1(_0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _1395_ (.A(_0733_),
    .B(_0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0741_));
 sky130_fd_sc_hd__and4_1 _1396_ (.A(net123),
    .B(_0739_),
    .C(_0740_),
    .D(_0741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _1397_ (.A1(net58),
    .A2(\tokenflow_inst.i6.ydata[74] ),
    .B1(\tokenflow_inst.i6.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0742_));
 sky130_fd_sc_hd__and3_1 _1398_ (.A(net58),
    .B(\tokenflow_inst.i6.ydata[22] ),
    .C(\tokenflow_inst.i6.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0743_));
 sky130_fd_sc_hd__inv_2 _1399_ (.A(_0743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0744_));
 sky130_fd_sc_hd__or2_1 _1400_ (.A(_0742_),
    .B(_0743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0745_));
 sky130_fd_sc_hd__a21oi_2 _1401_ (.A1(_0733_),
    .A2(_0738_),
    .B1(_0737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0746_));
 sky130_fd_sc_hd__a21o_1 _1402_ (.A1(_0740_),
    .A2(_0746_),
    .B1(_0745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0747_));
 sky130_fd_sc_hd__a31o_1 _1403_ (.A1(_0740_),
    .A2(_0745_),
    .A3(_0746_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0748_));
 sky130_fd_sc_hd__and2b_1 _1404_ (.A_N(_0748_),
    .B(_0747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__a21oi_1 _1405_ (.A1(net58),
    .A2(\tokenflow_inst.i6.ydata[75] ),
    .B1(\tokenflow_inst.i6.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0749_));
 sky130_fd_sc_hd__nand3_1 _1406_ (.A(net58),
    .B(\tokenflow_inst.i6.ydata[23] ),
    .C(\tokenflow_inst.i6.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2b_1 _1407_ (.A_N(_0749_),
    .B(_0750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0751_));
 sky130_fd_sc_hd__a21oi_1 _1408_ (.A1(_0744_),
    .A2(_0747_),
    .B1(_0751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0752_));
 sky130_fd_sc_hd__a31o_1 _1409_ (.A1(_0744_),
    .A2(_0747_),
    .A3(_0751_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_1 _1410_ (.A(_0752_),
    .B(_0753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0289_));
 sky130_fd_sc_hd__or2_1 _1411_ (.A(_0745_),
    .B(_0751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _1412_ (.A(_0740_),
    .B(_0754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0755_));
 sky130_fd_sc_hd__o221ai_2 _1413_ (.A1(_0744_),
    .A2(_0749_),
    .B1(_0754_),
    .B2(_0746_),
    .C1(_0750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0756_));
 sky130_fd_sc_hd__a21oi_1 _1414_ (.A1(net58),
    .A2(\tokenflow_inst.i6.ydata[76] ),
    .B1(\tokenflow_inst.i6.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0757_));
 sky130_fd_sc_hd__and3_1 _1415_ (.A(net58),
    .B(\tokenflow_inst.i6.ydata[76] ),
    .C(\tokenflow_inst.i6.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0758_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(_0758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0757_),
    .B(_0758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0760_));
 sky130_fd_sc_hd__or3_1 _1418_ (.A(_0755_),
    .B(_0756_),
    .C(_0760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0761_));
 sky130_fd_sc_hd__o21ai_1 _1419_ (.A1(_0755_),
    .A2(_0756_),
    .B1(_0760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0762_));
 sky130_fd_sc_hd__and3_1 _1420_ (.A(net104),
    .B(_0761_),
    .C(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_1 _1421_ (.A(net58),
    .B(\tokenflow_inst.i6.ydata[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0763_));
 sky130_fd_sc_hd__xor2_1 _1422_ (.A(\tokenflow_inst.i6.ydata[25] ),
    .B(_0763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0764_));
 sky130_fd_sc_hd__a21oi_1 _1423_ (.A1(_0759_),
    .A2(_0762_),
    .B1(_0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0765_));
 sky130_fd_sc_hd__a31o_1 _1424_ (.A1(_0759_),
    .A2(_0762_),
    .A3(_0764_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(_0765_),
    .B(_0766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0291_));
 sky130_fd_sc_hd__and2_1 _1426_ (.A(net117),
    .B(\tokenflow_inst.i6.ydata[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(net116),
    .B(\tokenflow_inst.i6.ydata[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__and2_1 _1428_ (.A(net145),
    .B(\tokenflow_inst.i6.ydata[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__and2_1 _1429_ (.A(net116),
    .B(\tokenflow_inst.i6.ydata[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__and2_1 _1430_ (.A(net145),
    .B(\tokenflow_inst.i6.ydata[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(net111),
    .B(\tokenflow_inst.i6.ydata[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__and2_1 _1432_ (.A(net112),
    .B(\tokenflow_inst.i6.ydata[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__and2_1 _1433_ (.A(net111),
    .B(\tokenflow_inst.i6.ydata[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _1434_ (.A(net110),
    .B(\tokenflow_inst.i6.ydata[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__and2_1 _1435_ (.A(net92),
    .B(\tokenflow_inst.i6.ydata[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _1436_ (.A(net96),
    .B(\tokenflow_inst.i6.ydata[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__and2_1 _1437_ (.A(net90),
    .B(\tokenflow_inst.i6.ydata[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__and2_1 _1438_ (.A(net90),
    .B(\tokenflow_inst.i6.ydata[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _1439_ (.A(net90),
    .B(\tokenflow_inst.i6.ydata[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__and2_1 _1440_ (.A(net90),
    .B(\tokenflow_inst.i6.ydata[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _1441_ (.A(net92),
    .B(\tokenflow_inst.i6.ydata[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__and2_1 _1442_ (.A(net92),
    .B(\tokenflow_inst.i6.ydata[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _1443_ (.A(net96),
    .B(\tokenflow_inst.i6.ydata[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _1444_ (.A(net97),
    .B(\tokenflow_inst.i6.ydata[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _1445_ (.A(net110),
    .B(\tokenflow_inst.i6.ydata[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__and2_1 _1446_ (.A(net97),
    .B(\tokenflow_inst.i6.ydata[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _1447_ (.A(net96),
    .B(\tokenflow_inst.i6.ydata[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _1448_ (.A(net96),
    .B(\tokenflow_inst.i6.ydata[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__and2_1 _1449_ (.A(net96),
    .B(\tokenflow_inst.i6.ydata[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__and2_1 _1450_ (.A(net93),
    .B(\tokenflow_inst.i6.ydata[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _1451_ (.A(net127),
    .B(\tokenflow_inst.i6.ydata[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _1452_ (.A(net129),
    .B(\tokenflow_inst.i6.ydata[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__and2_1 _1453_ (.A(net127),
    .B(\tokenflow_inst.i6.ydata[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _1454_ (.A(net125),
    .B(\tokenflow_inst.i6.ydata[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _1455_ (.A(net125),
    .B(\tokenflow_inst.i6.ydata[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__and2_1 _1456_ (.A(net122),
    .B(\tokenflow_inst.i6.ydata[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _1457_ (.A(net113),
    .B(\tokenflow_inst.i6.ydata[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _1458_ (.A(net114),
    .B(\tokenflow_inst.i6.ydata[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(net100),
    .B(\tokenflow_inst.i6.ydata[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _1460_ (.A(net100),
    .B(\tokenflow_inst.i6.ydata[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__and2_1 _1461_ (.A(net95),
    .B(\tokenflow_inst.i6.ydata[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _1462_ (.A(net103),
    .B(\tokenflow_inst.i6.ydata[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _1463_ (.A(net102),
    .B(\tokenflow_inst.i6.ydata[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__and2_1 _1464_ (.A(net102),
    .B(\tokenflow_inst.i6.ydata[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _1465_ (.A(net103),
    .B(\tokenflow_inst.i6.ydata[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _1466_ (.A(net104),
    .B(\tokenflow_inst.i6.ydata[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _1467_ (.A(net122),
    .B(\tokenflow_inst.i6.ydata[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _1468_ (.A(net123),
    .B(\tokenflow_inst.i6.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__and2_1 _1469_ (.A(net124),
    .B(\tokenflow_inst.i6.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__and2_1 _1470_ (.A(net128),
    .B(\tokenflow_inst.i6.ydata[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _1471_ (.A(net107),
    .B(\tokenflow_inst.i6.ydata[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _1472_ (.A(net107),
    .B(\tokenflow_inst.i6.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__and2_1 _1473_ (.A(net105),
    .B(\tokenflow_inst.i6.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _1474_ (.A(net105),
    .B(\tokenflow_inst.i6.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__and2_1 _1475_ (.A(net104),
    .B(\tokenflow_inst.i6.ydata[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__and2_1 _1476_ (.A(net129),
    .B(\tokenflow_inst.i3.ydata[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _1477_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _1478_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _1479_ (.A(net125),
    .B(\tokenflow_inst.i3.ydata[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _1480_ (.A(net125),
    .B(\tokenflow_inst.i3.ydata[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _1481_ (.A(net122),
    .B(\tokenflow_inst.i3.ydata[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _1482_ (.A(net122),
    .B(\tokenflow_inst.i3.ydata[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _1483_ (.A(net122),
    .B(\tokenflow_inst.i3.ydata[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _1484_ (.A(net100),
    .B(\tokenflow_inst.i3.ydata[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__and2_1 _1485_ (.A(net100),
    .B(\tokenflow_inst.i3.ydata[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _1486_ (.A(net102),
    .B(\tokenflow_inst.i3.ydata[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _1487_ (.A(net108),
    .B(\tokenflow_inst.i3.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _1488_ (.A(net102),
    .B(\tokenflow_inst.i3.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _1489_ (.A(net102),
    .B(\tokenflow_inst.i3.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0120_));
 sky130_fd_sc_hd__and2_1 _1490_ (.A(net106),
    .B(\tokenflow_inst.i3.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _1491_ (.A(net106),
    .B(\tokenflow_inst.i3.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _1492_ (.A(net122),
    .B(\tokenflow_inst.i3.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _1493_ (.A(net107),
    .B(\tokenflow_inst.i3.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _1494_ (.A(net124),
    .B(\tokenflow_inst.i3.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _1495_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0126_));
 sky130_fd_sc_hd__and2_1 _1496_ (.A(net124),
    .B(\tokenflow_inst.i3.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _1497_ (.A(net107),
    .B(\tokenflow_inst.i3.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _1498_ (.A(net106),
    .B(\tokenflow_inst.i3.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _1499_ (.A(net105),
    .B(\tokenflow_inst.i3.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__and2_1 _1500_ (.A(net104),
    .B(\tokenflow_inst.i3.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__and2_1 _1501_ (.A(net104),
    .B(\tokenflow_inst.i3.ydata[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _1502_ (.A(net117),
    .B(\tokenflow_inst.i3.ydata[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _1503_ (.A(net117),
    .B(\tokenflow_inst.i3.ydata[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _1504_ (.A(net116),
    .B(\tokenflow_inst.i3.ydata[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _1505_ (.A(net121),
    .B(\tokenflow_inst.i3.ydata[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _1506_ (.A(net115),
    .B(\tokenflow_inst.i3.ydata[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _1507_ (.A(net115),
    .B(\tokenflow_inst.i3.ydata[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__and2_1 _1508_ (.A(net111),
    .B(\tokenflow_inst.i3.ydata[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _1509_ (.A(net112),
    .B(\tokenflow_inst.i3.ydata[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__and2_1 _1510_ (.A(net111),
    .B(\tokenflow_inst.i3.ydata[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _1511_ (.A(net110),
    .B(\tokenflow_inst.i3.ydata[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _1512_ (.A(net92),
    .B(\tokenflow_inst.i3.ydata[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _1513_ (.A(net92),
    .B(\tokenflow_inst.i3.ydata[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__and2_1 _1514_ (.A(net90),
    .B(\tokenflow_inst.i3.ydata[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _1515_ (.A(net90),
    .B(\tokenflow_inst.i3.ydata[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _1516_ (.A(net90),
    .B(\tokenflow_inst.i3.ydata[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _1517_ (.A(net96),
    .B(\tokenflow_inst.i3.ydata[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _1518_ (.A(net92),
    .B(\tokenflow_inst.i3.ydata[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__and2_1 _1519_ (.A(net96),
    .B(\tokenflow_inst.i3.ydata[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _1520_ (.A(net96),
    .B(\tokenflow_inst.i3.ydata[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _1521_ (.A(net97),
    .B(\tokenflow_inst.i3.ydata[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _1522_ (.A(net110),
    .B(\tokenflow_inst.i3.ydata[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _1523_ (.A(net97),
    .B(\tokenflow_inst.i3.ydata[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _1524_ (.A(net98),
    .B(\tokenflow_inst.i3.ydata[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _1525_ (.A(net98),
    .B(\tokenflow_inst.i3.ydata[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _1526_ (.A(net98),
    .B(\tokenflow_inst.i3.ydata[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _1527_ (.A(net93),
    .B(\tokenflow_inst.i3.ydata[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__and2_1 _1528_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _1529_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__and2_1 _1530_ (.A(net127),
    .B(\tokenflow_inst.i3.ydata[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _1531_ (.A(net126),
    .B(\tokenflow_inst.i3.ydata[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _1532_ (.A(net126),
    .B(\tokenflow_inst.i3.ydata[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _1533_ (.A(net126),
    .B(\tokenflow_inst.i3.ydata[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _1534_ (.A(net120),
    .B(\tokenflow_inst.i3.ydata[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _1535_ (.A(net114),
    .B(\tokenflow_inst.i3.ydata[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _1536_ (.A(net130),
    .B(\tokenflow_inst.i3.ydata[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _1537_ (.A(net100),
    .B(\tokenflow_inst.i3.ydata[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _1538_ (.A(net101),
    .B(\tokenflow_inst.i3.ydata[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(net99),
    .B(\tokenflow_inst.i3.ydata[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _1540_ (.A(net102),
    .B(\tokenflow_inst.i3.ydata[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _1541_ (.A(net102),
    .B(\tokenflow_inst.i3.ydata[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _1542_ (.A(net103),
    .B(\tokenflow_inst.i3.ydata[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _1543_ (.A(net103),
    .B(\tokenflow_inst.i3.ydata[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _1544_ (.A(net108),
    .B(\tokenflow_inst.i3.ydata[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _1545_ (.A(net107),
    .B(\tokenflow_inst.i3.ydata[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(net124),
    .B(\tokenflow_inst.i3.ydata[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _1547_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__and2_1 _1548_ (.A(net128),
    .B(\tokenflow_inst.i3.ydata[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _1549_ (.A(net123),
    .B(\tokenflow_inst.i3.ydata[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _1550_ (.A(net106),
    .B(\tokenflow_inst.i3.ydata[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__and2_1 _1551_ (.A(net106),
    .B(\tokenflow_inst.i3.ydata[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__and2_1 _1552_ (.A(net104),
    .B(\tokenflow_inst.i3.ydata[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _1553_ (.A(net104),
    .B(\tokenflow_inst.i3.ydata[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__nor2_1 _1554_ (.A(net87),
    .B(\tokenflow_inst.i2.cg2.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0113_));
 sky130_fd_sc_hd__and2_4 _1555_ (.A(\tokenflow_inst.i78.cg_elem.q ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1556_ (.A(\tokenflow_inst.i78.d0_elem.inv_chain[3] ),
    .B(net119),
    .C(\tokenflow_inst.i78.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _1557_ (.A(net119),
    .B(\tokenflow_inst.i1.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _1558_ (.A1(\tokenflow_inst.i1.c.q ),
    .A2(net18),
    .B1(\tokenflow_inst.i2.cg1.q ),
    .B2(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_1 _1559_ (.A(net87),
    .B(\tokenflow_inst.i6.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0194_));
 sky130_fd_sc_hd__and2b_1 _1560_ (.A_N(\tokenflow_inst.i9.c.q ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_1 _1561_ (.A(net86),
    .B(\tokenflow_inst.i1.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0033_));
 sky130_fd_sc_hd__and2_4 _1562_ (.A(\tokenflow_inst.i2.cg2.a ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and2_1 _1563_ (.A(net126),
    .B(\tokenflow_inst.i11.i.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1564_ (.A(net126),
    .B(\tokenflow_inst.i11.i.d0.inv_chain[1] ),
    .C(\tokenflow_inst.i11.i.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _1565_ (.A(net119),
    .B(\tokenflow_inst.ii3.i.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1566_ (.A(net119),
    .B(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ),
    .C(\tokenflow_inst.ii3.i.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__nor2_1 _1567_ (.A(net86),
    .B(\tokenflow_inst.ii3.i.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0380_));
 sky130_fd_sc_hd__and2_1 _1568_ (.A(net118),
    .B(\tokenflow_inst.ii1.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1569_ (.A(net118),
    .B(\tokenflow_inst.ii1.d0_elem.inv_chain[2] ),
    .C(\tokenflow_inst.ii1.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _1570_ (.A(net118),
    .B(\tokenflow_inst.ii2.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(net86),
    .B(\tokenflow_inst.ii1.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0352_));
 sky130_fd_sc_hd__xor2_4 _1572_ (.A(\tokenflow_inst.i3.ydata[0] ),
    .B(\tokenflow_inst.i3.ydata[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__xor2_4 _1573_ (.A(\tokenflow_inst.i3.ydata[1] ),
    .B(\tokenflow_inst.i3.ydata[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__xor2_4 _1574_ (.A(\tokenflow_inst.i3.ydata[2] ),
    .B(\tokenflow_inst.i3.ydata[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__xor2_4 _1575_ (.A(\tokenflow_inst.i3.ydata[3] ),
    .B(\tokenflow_inst.i3.ydata[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__xor2_4 _1576_ (.A(\tokenflow_inst.i3.ydata[4] ),
    .B(\tokenflow_inst.i3.ydata[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__xor2_4 _1577_ (.A(\tokenflow_inst.i3.ydata[5] ),
    .B(\tokenflow_inst.i3.ydata[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__xor2_4 _1578_ (.A(\tokenflow_inst.i3.ydata[6] ),
    .B(\tokenflow_inst.i3.ydata[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__xor2_4 _1579_ (.A(\tokenflow_inst.i3.ydata[7] ),
    .B(\tokenflow_inst.i3.ydata[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__xor2_4 _1580_ (.A(\tokenflow_inst.i3.ydata[8] ),
    .B(\tokenflow_inst.i3.ydata[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__xor2_4 _1581_ (.A(\tokenflow_inst.i3.ydata[9] ),
    .B(\tokenflow_inst.i3.ydata[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__xor2_4 _1582_ (.A(\tokenflow_inst.i3.ydata[10] ),
    .B(\tokenflow_inst.i3.ydata[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__or4_1 _1583_ (.A(\tokenflow_inst.i3.ydata[48] ),
    .B(\tokenflow_inst.i3.ydata[49] ),
    .C(\tokenflow_inst.i3.ydata[50] ),
    .D(\tokenflow_inst.i3.ydata[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0767_));
 sky130_fd_sc_hd__or4_1 _1584_ (.A(\tokenflow_inst.i3.ydata[44] ),
    .B(\tokenflow_inst.i3.ydata[45] ),
    .C(\tokenflow_inst.i3.ydata[46] ),
    .D(\tokenflow_inst.i3.ydata[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0768_));
 sky130_fd_sc_hd__or4_1 _1585_ (.A(\tokenflow_inst.i3.ydata[40] ),
    .B(\tokenflow_inst.i3.ydata[41] ),
    .C(\tokenflow_inst.i3.ydata[42] ),
    .D(\tokenflow_inst.i3.ydata[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0769_));
 sky130_fd_sc_hd__or3_1 _1586_ (.A(_0767_),
    .B(_0768_),
    .C(_0769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0770_));
 sky130_fd_sc_hd__or4_1 _1587_ (.A(\tokenflow_inst.i3.ydata[28] ),
    .B(\tokenflow_inst.i3.ydata[29] ),
    .C(\tokenflow_inst.i3.ydata[30] ),
    .D(\tokenflow_inst.i3.ydata[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0771_));
 sky130_fd_sc_hd__or4_1 _1588_ (.A(\tokenflow_inst.i3.ydata[36] ),
    .B(\tokenflow_inst.i3.ydata[37] ),
    .C(\tokenflow_inst.i3.ydata[38] ),
    .D(\tokenflow_inst.i3.ydata[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0772_));
 sky130_fd_sc_hd__or4_1 _1589_ (.A(\tokenflow_inst.i3.ydata[32] ),
    .B(\tokenflow_inst.i3.ydata[33] ),
    .C(\tokenflow_inst.i3.ydata[34] ),
    .D(\tokenflow_inst.i3.ydata[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0773_));
 sky130_fd_sc_hd__or4_1 _1590_ (.A(\tokenflow_inst.i3.ydata[26] ),
    .B(\tokenflow_inst.i3.ydata[27] ),
    .C(_0771_),
    .D(_0772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0774_));
 sky130_fd_sc_hd__nor3_1 _1591_ (.A(_0770_),
    .B(_0773_),
    .C(_0774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0775_));
 sky130_fd_sc_hd__and3_1 _1592_ (.A(\tokenflow_inst.i3.d0_elem.inv_chain[3] ),
    .B(\tokenflow_inst.i2.cg2.a ),
    .C(_0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i10.cg.b ));
 sky130_fd_sc_hd__and2_1 _1593_ (.A(net125),
    .B(\tokenflow_inst.i10.cg.b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _1594_ (.A(net86),
    .B(\tokenflow_inst.i11.i.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0028_));
 sky130_fd_sc_hd__and2_1 _1595_ (.A(net126),
    .B(\tokenflow_inst.i10.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i10.d0.inv_chain[0] ));
 sky130_fd_sc_hd__and2_1 _1596_ (.A(net128),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_1 _1597_ (.A(net87),
    .B(\tokenflow_inst.i78.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0271_));
 sky130_fd_sc_hd__and2_4 _1598_ (.A(net115),
    .B(\tokenflow_inst.i8.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1599_ (.A(\tokenflow_inst.i8.d0_elem.inv_chain[52] ),
    .B(net118),
    .C(\tokenflow_inst.i8.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__nor2_1 _1600_ (.A(net87),
    .B(\tokenflow_inst.i2.cg2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0272_));
 sky130_fd_sc_hd__nor2_1 _1601_ (.A(net86),
    .B(\tokenflow_inst.i8.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0195_));
 sky130_fd_sc_hd__and2_1 _1602_ (.A(net115),
    .B(\tokenflow_inst.i6.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[0] ));
 sky130_fd_sc_hd__and3_1 _1603_ (.A(net115),
    .B(\tokenflow_inst.i6.cg_elem.q ),
    .C(\tokenflow_inst.i6.d0_elem.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__and3b_1 _1604_ (.A_N(_0775_),
    .B(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .C(\tokenflow_inst.i3.d0_elem.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__dlxtn_1 _1605_ (.D(_0062_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[34] ));
 sky130_fd_sc_hd__dlxtn_1 _1606_ (.D(_0063_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[35] ));
 sky130_fd_sc_hd__dlxtn_1 _1607_ (.D(_0064_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[36] ));
 sky130_fd_sc_hd__dlxtn_1 _1608_ (.D(_0065_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[37] ));
 sky130_fd_sc_hd__dlxtn_1 _1609_ (.D(_0066_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[38] ));
 sky130_fd_sc_hd__dlxtn_1 _1610_ (.D(_0067_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[39] ));
 sky130_fd_sc_hd__dlxtn_1 _1611_ (.D(_0069_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[40] ));
 sky130_fd_sc_hd__dlxtn_1 _1612_ (.D(_0070_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[41] ));
 sky130_fd_sc_hd__dlxtn_1 _1613_ (.D(_0071_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[42] ));
 sky130_fd_sc_hd__dlxtn_1 _1614_ (.D(_0072_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[43] ));
 sky130_fd_sc_hd__dlxtn_1 _1615_ (.D(_0073_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[44] ));
 sky130_fd_sc_hd__dlxtn_1 _1616_ (.D(_0074_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[45] ));
 sky130_fd_sc_hd__dlxtn_1 _1617_ (.D(_0075_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[46] ));
 sky130_fd_sc_hd__dlxtn_1 _1618_ (.D(_0076_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[47] ));
 sky130_fd_sc_hd__dlxtn_1 _1619_ (.D(_0077_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[48] ));
 sky130_fd_sc_hd__dlxtn_1 _1620_ (.D(_0078_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[49] ));
 sky130_fd_sc_hd__dlxtn_1 _1621_ (.D(_0080_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[50] ));
 sky130_fd_sc_hd__dlxtn_1 _1622_ (.D(_0081_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[51] ));
 sky130_fd_sc_hd__dlxtn_1 _1623_ (.D(_0082_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[52] ));
 sky130_fd_sc_hd__dlxtn_1 _1624_ (.D(_0083_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[53] ));
 sky130_fd_sc_hd__dlxtn_1 _1625_ (.D(_0084_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[54] ));
 sky130_fd_sc_hd__dlxtn_1 _1626_ (.D(_0085_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[55] ));
 sky130_fd_sc_hd__dlxtn_1 _1627_ (.D(_0086_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[56] ));
 sky130_fd_sc_hd__dlxtn_1 _1628_ (.D(_0087_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[57] ));
 sky130_fd_sc_hd__dlxtn_1 _1629_ (.D(_0088_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[58] ));
 sky130_fd_sc_hd__dlxtn_1 _1630_ (.D(_0089_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[59] ));
 sky130_fd_sc_hd__dlxtn_1 _1631_ (.D(_0091_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[60] ));
 sky130_fd_sc_hd__dlxtn_1 _1632_ (.D(_0092_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[61] ));
 sky130_fd_sc_hd__dlxtn_1 _1633_ (.D(_0093_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[62] ));
 sky130_fd_sc_hd__dlxtn_1 _1634_ (.D(_0094_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[63] ));
 sky130_fd_sc_hd__dlxtn_1 _1635_ (.D(_0095_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[64] ));
 sky130_fd_sc_hd__dlxtn_1 _1636_ (.D(_0096_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[65] ));
 sky130_fd_sc_hd__dlxtn_1 _1637_ (.D(_0097_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[66] ));
 sky130_fd_sc_hd__dlxtn_1 _1638_ (.D(_0098_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[67] ));
 sky130_fd_sc_hd__dlxtn_1 _1639_ (.D(_0099_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[68] ));
 sky130_fd_sc_hd__dlxtn_1 _1640_ (.D(_0100_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[69] ));
 sky130_fd_sc_hd__dlxtn_1 _1641_ (.D(_0102_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[70] ));
 sky130_fd_sc_hd__dlxtn_1 _1642_ (.D(_0103_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[71] ));
 sky130_fd_sc_hd__dlxtn_1 _1643_ (.D(_0104_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[72] ));
 sky130_fd_sc_hd__dlxtn_1 _1644_ (.D(_0105_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[73] ));
 sky130_fd_sc_hd__dlxtn_1 _1645_ (.D(_0106_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[74] ));
 sky130_fd_sc_hd__dlxtn_1 _1646_ (.D(_0107_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[75] ));
 sky130_fd_sc_hd__dlxtn_1 _1647_ (.D(_0108_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[76] ));
 sky130_fd_sc_hd__dlxtn_1 _1648_ (.D(_0109_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[77] ));
 sky130_fd_sc_hd__dlxtn_1 _1649_ (.D(_0382_),
    .GATE_N(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1650_ (.D(_0393_),
    .GATE_N(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_2 _1651_ (.D(_0400_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1652_ (.D(_0401_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_2 _1653_ (.D(_0402_),
    .GATE_N(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1654_ (.D(_0403_),
    .GATE_N(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1655_ (.D(_0404_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1656_ (.D(_0405_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1657_ (.D(_0406_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1658_ (.D(_0407_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1659_ (.D(_0383_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1660_ (.D(_0384_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1661_ (.D(_0385_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_2 _1662_ (.D(_0386_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_2 _1663_ (.D(_0387_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1664_ (.D(_0388_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_2 _1665_ (.D(_0389_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1666_ (.D(_0390_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_2 _1667_ (.D(_0391_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1668_ (.D(_0392_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_2 _1669_ (.D(_0394_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1670_ (.D(_0395_),
    .GATE_N(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1671_ (.D(_0396_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_2 _1672_ (.D(_0397_),
    .GATE_N(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1673_ (.D(_0398_),
    .GATE_N(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1674_ (.D(_0399_),
    .GATE_N(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii3.i.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1675_ (.D(_0354_),
    .GATE_N(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1676_ (.D(_0365_),
    .GATE_N(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_1 _1677_ (.D(_0372_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1678_ (.D(_0373_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1679_ (.D(_0374_),
    .GATE_N(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1680_ (.D(_0375_),
    .GATE_N(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1681_ (.D(_0376_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1682_ (.D(_0377_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1683_ (.D(_0378_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1684_ (.D(_0379_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1685_ (.D(_0355_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1686_ (.D(_0356_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1687_ (.D(_0357_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1688_ (.D(_0358_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1689_ (.D(_0359_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1690_ (.D(_0360_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1691_ (.D(_0361_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1692_ (.D(_0362_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1693_ (.D(_0363_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1694_ (.D(_0364_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1695_ (.D(_0366_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1696_ (.D(_0367_),
    .GATE_N(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1697_ (.D(_0368_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1698_ (.D(_0369_),
    .GATE_N(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1699_ (.D(_0370_),
    .GATE_N(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1700_ (.D(_0371_),
    .GATE_N(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii2.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1701_ (.D(_0000_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1702_ (.D(_0011_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_1 _1703_ (.D(_0018_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1704_ (.D(_0019_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1705_ (.D(_0020_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1706_ (.D(_0021_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1707_ (.D(_0022_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1708_ (.D(_0023_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1709_ (.D(_0024_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1710_ (.D(_0025_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1711_ (.D(_0001_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1712_ (.D(_0002_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1713_ (.D(_0003_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1714_ (.D(_0004_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1715_ (.D(_0005_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1716_ (.D(_0006_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1717_ (.D(_0007_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1718_ (.D(_0008_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1719_ (.D(_0009_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1720_ (.D(_0010_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1721_ (.D(_0012_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1722_ (.D(_0013_),
    .GATE_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1723_ (.D(_0014_),
    .GATE_N(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1724_ (.D(_0015_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1725_ (.D(_0016_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1726_ (.D(_0017_),
    .GATE_N(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.ii1.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1727_ (.D(_0274_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1728_ (.D(_0285_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_1 _1729_ (.D(_0296_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1730_ (.D(_0307_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1731_ (.D(_0318_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1732_ (.D(_0327_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1733_ (.D(_0338_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1734_ (.D(_0347_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1735_ (.D(_0348_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1736_ (.D(_0349_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1737_ (.D(_0275_),
    .GATE_N(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1738_ (.D(_0276_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1739_ (.D(_0277_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1740_ (.D(_0278_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1741_ (.D(_0279_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1742_ (.D(_0280_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1743_ (.D(_0281_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1744_ (.D(_0282_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1745_ (.D(_0283_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1746_ (.D(_0284_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1747_ (.D(_0286_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1748_ (.D(_0287_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1749_ (.D(_0288_),
    .GATE_N(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1750_ (.D(_0289_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1751_ (.D(_0290_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1752_ (.D(_0291_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1753_ (.D(_0292_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[26] ));
 sky130_fd_sc_hd__dlxtn_1 _1754_ (.D(_0293_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[27] ));
 sky130_fd_sc_hd__dlxtn_1 _1755_ (.D(_0294_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[28] ));
 sky130_fd_sc_hd__dlxtn_1 _1756_ (.D(_0295_),
    .GATE_N(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[29] ));
 sky130_fd_sc_hd__dlxtn_1 _1757_ (.D(_0297_),
    .GATE_N(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[30] ));
 sky130_fd_sc_hd__dlxtn_1 _1758_ (.D(_0298_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[31] ));
 sky130_fd_sc_hd__dlxtn_1 _1759_ (.D(_0299_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[32] ));
 sky130_fd_sc_hd__dlxtn_1 _1760_ (.D(_0300_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[33] ));
 sky130_fd_sc_hd__dlxtn_1 _1761_ (.D(_0301_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[34] ));
 sky130_fd_sc_hd__dlxtn_1 _1762_ (.D(_0302_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[35] ));
 sky130_fd_sc_hd__dlxtn_1 _1763_ (.D(_0303_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[36] ));
 sky130_fd_sc_hd__dlxtn_1 _1764_ (.D(_0304_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[37] ));
 sky130_fd_sc_hd__dlxtn_1 _1765_ (.D(_0305_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[38] ));
 sky130_fd_sc_hd__dlxtn_1 _1766_ (.D(_0306_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[39] ));
 sky130_fd_sc_hd__dlxtn_1 _1767_ (.D(_0308_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[40] ));
 sky130_fd_sc_hd__dlxtn_1 _1768_ (.D(_0309_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[41] ));
 sky130_fd_sc_hd__dlxtn_1 _1769_ (.D(_0310_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[42] ));
 sky130_fd_sc_hd__dlxtn_1 _1770_ (.D(_0311_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[43] ));
 sky130_fd_sc_hd__dlxtn_1 _1771_ (.D(_0312_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[44] ));
 sky130_fd_sc_hd__dlxtn_1 _1772_ (.D(_0313_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[45] ));
 sky130_fd_sc_hd__dlxtn_1 _1773_ (.D(_0314_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[46] ));
 sky130_fd_sc_hd__dlxtn_1 _1774_ (.D(_0315_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[47] ));
 sky130_fd_sc_hd__dlxtn_1 _1775_ (.D(_0316_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[48] ));
 sky130_fd_sc_hd__dlxtn_1 _1776_ (.D(_0317_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[49] ));
 sky130_fd_sc_hd__dlxtn_1 _1777_ (.D(_0319_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[50] ));
 sky130_fd_sc_hd__dlxtn_1 _1778_ (.D(_0320_),
    .GATE_N(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[53] ));
 sky130_fd_sc_hd__dlxtn_1 _1779_ (.D(_0321_),
    .GATE_N(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[54] ));
 sky130_fd_sc_hd__dlxtn_1 _1780_ (.D(_0322_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[55] ));
 sky130_fd_sc_hd__dlxtn_1 _1781_ (.D(_0323_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[56] ));
 sky130_fd_sc_hd__dlxtn_1 _1782_ (.D(_0324_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[57] ));
 sky130_fd_sc_hd__dlxtn_1 _1783_ (.D(_0325_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[58] ));
 sky130_fd_sc_hd__dlxtn_1 _1784_ (.D(_0326_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[59] ));
 sky130_fd_sc_hd__dlxtn_1 _1785_ (.D(_0328_),
    .GATE_N(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[60] ));
 sky130_fd_sc_hd__dlxtn_1 _1786_ (.D(_0329_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[61] ));
 sky130_fd_sc_hd__dlxtn_1 _1787_ (.D(_0330_),
    .GATE_N(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[62] ));
 sky130_fd_sc_hd__dlxtn_1 _1788_ (.D(_0331_),
    .GATE_N(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[63] ));
 sky130_fd_sc_hd__dlxtn_1 _1789_ (.D(_0332_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[64] ));
 sky130_fd_sc_hd__dlxtn_1 _1790_ (.D(_0333_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[65] ));
 sky130_fd_sc_hd__dlxtn_1 _1791_ (.D(_0334_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[66] ));
 sky130_fd_sc_hd__dlxtn_1 _1792_ (.D(_0335_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[67] ));
 sky130_fd_sc_hd__dlxtn_1 _1793_ (.D(_0336_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[68] ));
 sky130_fd_sc_hd__dlxtn_1 _1794_ (.D(_0337_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[69] ));
 sky130_fd_sc_hd__dlxtn_1 _1795_ (.D(_0339_),
    .GATE_N(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[70] ));
 sky130_fd_sc_hd__dlxtn_1 _1796_ (.D(_0340_),
    .GATE_N(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[71] ));
 sky130_fd_sc_hd__dlxtn_1 _1797_ (.D(_0341_),
    .GATE_N(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[72] ));
 sky130_fd_sc_hd__dlxtn_1 _1798_ (.D(_0342_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[73] ));
 sky130_fd_sc_hd__dlxtn_1 _1799_ (.D(_0343_),
    .GATE_N(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[74] ));
 sky130_fd_sc_hd__dlxtn_1 _1800_ (.D(_0344_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[75] ));
 sky130_fd_sc_hd__dlxtn_1 _1801_ (.D(_0345_),
    .GATE_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[76] ));
 sky130_fd_sc_hd__dlxtn_1 _1802_ (.D(_0346_),
    .GATE_N(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i8.ydata[77] ));
 sky130_fd_sc_hd__dlxtn_1 _1803_ (.D(_0197_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1804_ (.D(_0208_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_1 _1805_ (.D(_0219_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1806_ (.D(_0230_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1807_ (.D(_0241_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1808_ (.D(_0248_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1809_ (.D(_0259_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1810_ (.D(_0268_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1811_ (.D(_0269_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1812_ (.D(_0270_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1813_ (.D(_0198_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1814_ (.D(_0199_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1815_ (.D(_0200_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1816_ (.D(_0201_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1817_ (.D(_0202_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1818_ (.D(_0203_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1819_ (.D(_0204_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1820_ (.D(_0205_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1821_ (.D(_0206_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1822_ (.D(_0207_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1823_ (.D(_0209_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1824_ (.D(_0210_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1825_ (.D(_0211_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1826_ (.D(_0212_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1827_ (.D(_0213_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1828_ (.D(_0214_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1829_ (.D(_0215_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[26] ));
 sky130_fd_sc_hd__dlxtn_1 _1830_ (.D(_0216_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[27] ));
 sky130_fd_sc_hd__dlxtn_1 _1831_ (.D(_0217_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[28] ));
 sky130_fd_sc_hd__dlxtn_1 _1832_ (.D(_0218_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[29] ));
 sky130_fd_sc_hd__dlxtn_1 _1833_ (.D(_0220_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[30] ));
 sky130_fd_sc_hd__dlxtn_1 _1834_ (.D(_0221_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[31] ));
 sky130_fd_sc_hd__dlxtn_1 _1835_ (.D(_0222_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[32] ));
 sky130_fd_sc_hd__dlxtn_1 _1836_ (.D(_0223_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[33] ));
 sky130_fd_sc_hd__dlxtn_1 _1837_ (.D(_0224_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[34] ));
 sky130_fd_sc_hd__dlxtn_1 _1838_ (.D(_0225_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[35] ));
 sky130_fd_sc_hd__dlxtn_1 _1839_ (.D(_0226_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[36] ));
 sky130_fd_sc_hd__dlxtn_1 _1840_ (.D(_0227_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[37] ));
 sky130_fd_sc_hd__dlxtn_1 _1841_ (.D(_0228_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[38] ));
 sky130_fd_sc_hd__dlxtn_1 _1842_ (.D(_0229_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[39] ));
 sky130_fd_sc_hd__dlxtn_1 _1843_ (.D(_0231_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[40] ));
 sky130_fd_sc_hd__dlxtn_1 _1844_ (.D(_0232_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[41] ));
 sky130_fd_sc_hd__dlxtn_1 _1845_ (.D(_0233_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[42] ));
 sky130_fd_sc_hd__dlxtn_1 _1846_ (.D(_0234_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[43] ));
 sky130_fd_sc_hd__dlxtn_1 _1847_ (.D(_0235_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[44] ));
 sky130_fd_sc_hd__dlxtn_1 _1848_ (.D(_0236_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[45] ));
 sky130_fd_sc_hd__dlxtn_1 _1849_ (.D(_0237_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[46] ));
 sky130_fd_sc_hd__dlxtn_1 _1850_ (.D(_0238_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[47] ));
 sky130_fd_sc_hd__dlxtn_1 _1851_ (.D(_0239_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[48] ));
 sky130_fd_sc_hd__dlxtn_1 _1852_ (.D(_0240_),
    .GATE_N(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[49] ));
 sky130_fd_sc_hd__dlxtn_1 _1853_ (.D(_0242_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[54] ));
 sky130_fd_sc_hd__dlxtn_1 _1854_ (.D(_0243_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[55] ));
 sky130_fd_sc_hd__dlxtn_1 _1855_ (.D(_0244_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[56] ));
 sky130_fd_sc_hd__dlxtn_1 _1856_ (.D(_0245_),
    .GATE_N(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[57] ));
 sky130_fd_sc_hd__dlxtn_1 _1857_ (.D(_0246_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[58] ));
 sky130_fd_sc_hd__dlxtn_1 _1858_ (.D(_0247_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[59] ));
 sky130_fd_sc_hd__dlxtn_1 _1859_ (.D(_0249_),
    .GATE_N(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[60] ));
 sky130_fd_sc_hd__dlxtn_1 _1860_ (.D(_0250_),
    .GATE_N(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[61] ));
 sky130_fd_sc_hd__dlxtn_1 _1861_ (.D(_0251_),
    .GATE_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[62] ));
 sky130_fd_sc_hd__dlxtn_1 _1862_ (.D(_0252_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[63] ));
 sky130_fd_sc_hd__dlxtn_1 _1863_ (.D(_0253_),
    .GATE_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[64] ));
 sky130_fd_sc_hd__dlxtn_1 _1864_ (.D(_0254_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[65] ));
 sky130_fd_sc_hd__dlxtn_1 _1865_ (.D(_0255_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[66] ));
 sky130_fd_sc_hd__dlxtn_1 _1866_ (.D(_0256_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[67] ));
 sky130_fd_sc_hd__dlxtn_1 _1867_ (.D(_0257_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[68] ));
 sky130_fd_sc_hd__dlxtn_1 _1868_ (.D(_0258_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[69] ));
 sky130_fd_sc_hd__dlxtn_1 _1869_ (.D(_0260_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[70] ));
 sky130_fd_sc_hd__dlxtn_1 _1870_ (.D(_0261_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[71] ));
 sky130_fd_sc_hd__dlxtn_1 _1871_ (.D(_0262_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[72] ));
 sky130_fd_sc_hd__dlxtn_1 _1872_ (.D(_0263_),
    .GATE_N(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[73] ));
 sky130_fd_sc_hd__dlxtn_1 _1873_ (.D(_0264_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[74] ));
 sky130_fd_sc_hd__dlxtn_1 _1874_ (.D(_0265_),
    .GATE_N(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[75] ));
 sky130_fd_sc_hd__dlxtn_1 _1875_ (.D(_0266_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[76] ));
 sky130_fd_sc_hd__dlxtn_1 _1876_ (.D(_0267_),
    .GATE_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i78.ydata[77] ));
 sky130_fd_sc_hd__dlxtn_1 _1877_ (.D(_0116_),
    .GATE_N(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_1 _1878_ (.D(_0127_),
    .GATE_N(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_1 _1879_ (.D(_0138_),
    .GATE_N(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1880_ (.D(_0149_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1881_ (.D(_0160_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_1 _1882_ (.D(_0171_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_1 _1883_ (.D(_0182_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_1 _1884_ (.D(_0191_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_1 _1885_ (.D(_0192_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_1 _1886_ (.D(_0193_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_1 _1887_ (.D(_0117_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1888_ (.D(_0118_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1889_ (.D(_0119_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1890_ (.D(_0120_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1891_ (.D(_0121_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1892_ (.D(_0122_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1893_ (.D(_0123_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1894_ (.D(_0124_),
    .GATE_N(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1895_ (.D(_0125_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1896_ (.D(_0126_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1897_ (.D(_0128_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1898_ (.D(_0129_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1899_ (.D(_0130_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1900_ (.D(_0131_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1901_ (.D(_0132_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1902_ (.D(_0133_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1903_ (.D(_0134_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[26] ));
 sky130_fd_sc_hd__dlxtn_1 _1904_ (.D(_0135_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[27] ));
 sky130_fd_sc_hd__dlxtn_1 _1905_ (.D(_0136_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[28] ));
 sky130_fd_sc_hd__dlxtn_1 _1906_ (.D(_0137_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[29] ));
 sky130_fd_sc_hd__dlxtn_1 _1907_ (.D(_0139_),
    .GATE_N(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[30] ));
 sky130_fd_sc_hd__dlxtn_1 _1908_ (.D(_0140_),
    .GATE_N(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[31] ));
 sky130_fd_sc_hd__dlxtn_1 _1909_ (.D(_0141_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[32] ));
 sky130_fd_sc_hd__dlxtn_1 _1910_ (.D(_0142_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[33] ));
 sky130_fd_sc_hd__dlxtn_1 _1911_ (.D(_0143_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[34] ));
 sky130_fd_sc_hd__dlxtn_1 _1912_ (.D(_0144_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[35] ));
 sky130_fd_sc_hd__dlxtn_1 _1913_ (.D(_0145_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[36] ));
 sky130_fd_sc_hd__dlxtn_1 _1914_ (.D(_0146_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[37] ));
 sky130_fd_sc_hd__dlxtn_1 _1915_ (.D(_0147_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[38] ));
 sky130_fd_sc_hd__dlxtn_1 _1916_ (.D(_0148_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[39] ));
 sky130_fd_sc_hd__dlxtn_1 _1917_ (.D(_0150_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[40] ));
 sky130_fd_sc_hd__dlxtn_1 _1918_ (.D(_0151_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[41] ));
 sky130_fd_sc_hd__dlxtn_1 _1919_ (.D(_0152_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[42] ));
 sky130_fd_sc_hd__dlxtn_1 _1920_ (.D(_0153_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[43] ));
 sky130_fd_sc_hd__dlxtn_1 _1921_ (.D(_0154_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[44] ));
 sky130_fd_sc_hd__dlxtn_1 _1922_ (.D(_0155_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[45] ));
 sky130_fd_sc_hd__dlxtn_1 _1923_ (.D(_0156_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[46] ));
 sky130_fd_sc_hd__dlxtn_1 _1924_ (.D(_0157_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[47] ));
 sky130_fd_sc_hd__dlxtn_1 _1925_ (.D(_0158_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[48] ));
 sky130_fd_sc_hd__dlxtn_1 _1926_ (.D(_0159_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[49] ));
 sky130_fd_sc_hd__dlxtn_1 _1927_ (.D(_0161_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[50] ));
 sky130_fd_sc_hd__dlxtn_1 _1928_ (.D(_0162_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[51] ));
 sky130_fd_sc_hd__dlxtn_1 _1929_ (.D(_0163_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[52] ));
 sky130_fd_sc_hd__dlxtn_1 _1930_ (.D(_0164_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[53] ));
 sky130_fd_sc_hd__dlxtn_1 _1931_ (.D(_0165_),
    .GATE_N(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[54] ));
 sky130_fd_sc_hd__dlxtn_1 _1932_ (.D(_0166_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[55] ));
 sky130_fd_sc_hd__dlxtn_1 _1933_ (.D(_0167_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[56] ));
 sky130_fd_sc_hd__dlxtn_1 _1934_ (.D(_0168_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[57] ));
 sky130_fd_sc_hd__dlxtn_1 _1935_ (.D(_0169_),
    .GATE_N(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[58] ));
 sky130_fd_sc_hd__dlxtn_1 _1936_ (.D(_0170_),
    .GATE_N(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[59] ));
 sky130_fd_sc_hd__dlxtn_1 _1937_ (.D(_0172_),
    .GATE_N(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[60] ));
 sky130_fd_sc_hd__dlxtn_1 _1938_ (.D(_0173_),
    .GATE_N(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[61] ));
 sky130_fd_sc_hd__dlxtn_1 _1939_ (.D(_0174_),
    .GATE_N(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[62] ));
 sky130_fd_sc_hd__dlxtn_1 _1940_ (.D(_0175_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[63] ));
 sky130_fd_sc_hd__dlxtn_1 _1941_ (.D(_0176_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[64] ));
 sky130_fd_sc_hd__dlxtn_1 _1942_ (.D(_0177_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[65] ));
 sky130_fd_sc_hd__dlxtn_1 _1943_ (.D(_0178_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[66] ));
 sky130_fd_sc_hd__dlxtn_1 _1944_ (.D(_0179_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[67] ));
 sky130_fd_sc_hd__dlxtn_1 _1945_ (.D(_0180_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[68] ));
 sky130_fd_sc_hd__dlxtn_1 _1946_ (.D(_0181_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[69] ));
 sky130_fd_sc_hd__dlxtn_1 _1947_ (.D(_0183_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[70] ));
 sky130_fd_sc_hd__dlxtn_1 _1948_ (.D(_0184_),
    .GATE_N(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[71] ));
 sky130_fd_sc_hd__dlxtn_1 _1949_ (.D(_0185_),
    .GATE_N(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[72] ));
 sky130_fd_sc_hd__dlxtn_1 _1950_ (.D(_0186_),
    .GATE_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[73] ));
 sky130_fd_sc_hd__dlxtn_1 _1951_ (.D(_0187_),
    .GATE_N(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[74] ));
 sky130_fd_sc_hd__dlxtn_1 _1952_ (.D(_0188_),
    .GATE_N(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[75] ));
 sky130_fd_sc_hd__dlxtn_1 _1953_ (.D(_0189_),
    .GATE_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[76] ));
 sky130_fd_sc_hd__dlxtn_1 _1954_ (.D(_0190_),
    .GATE_N(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i6.ydata[77] ));
 sky130_fd_sc_hd__dlxtn_2 _1955_ (.D(_0035_),
    .GATE_N(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[0] ));
 sky130_fd_sc_hd__dlxtn_2 _1956_ (.D(_0046_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[1] ));
 sky130_fd_sc_hd__dlxtn_2 _1957_ (.D(_0057_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[2] ));
 sky130_fd_sc_hd__dlxtn_1 _1958_ (.D(_0068_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[3] ));
 sky130_fd_sc_hd__dlxtn_1 _1959_ (.D(_0079_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[4] ));
 sky130_fd_sc_hd__dlxtn_2 _1960_ (.D(_0090_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[5] ));
 sky130_fd_sc_hd__dlxtn_2 _1961_ (.D(_0101_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[6] ));
 sky130_fd_sc_hd__dlxtn_2 _1962_ (.D(_0110_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[7] ));
 sky130_fd_sc_hd__dlxtn_2 _1963_ (.D(_0111_),
    .GATE_N(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[8] ));
 sky130_fd_sc_hd__dlxtn_2 _1964_ (.D(_0112_),
    .GATE_N(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[9] ));
 sky130_fd_sc_hd__dlxtn_2 _1965_ (.D(_0036_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[10] ));
 sky130_fd_sc_hd__dlxtn_1 _1966_ (.D(_0037_),
    .GATE_N(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[11] ));
 sky130_fd_sc_hd__dlxtn_1 _1967_ (.D(_0038_),
    .GATE_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[12] ));
 sky130_fd_sc_hd__dlxtn_1 _1968_ (.D(_0039_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[13] ));
 sky130_fd_sc_hd__dlxtn_1 _1969_ (.D(_0040_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[14] ));
 sky130_fd_sc_hd__dlxtn_1 _1970_ (.D(_0041_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[15] ));
 sky130_fd_sc_hd__dlxtn_1 _1971_ (.D(_0042_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[16] ));
 sky130_fd_sc_hd__dlxtn_1 _1972_ (.D(_0043_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[17] ));
 sky130_fd_sc_hd__dlxtn_1 _1973_ (.D(_0044_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[18] ));
 sky130_fd_sc_hd__dlxtn_1 _1974_ (.D(_0045_),
    .GATE_N(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[19] ));
 sky130_fd_sc_hd__dlxtn_1 _1975_ (.D(_0047_),
    .GATE_N(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[20] ));
 sky130_fd_sc_hd__dlxtn_1 _1976_ (.D(_0048_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[21] ));
 sky130_fd_sc_hd__dlxtn_1 _1977_ (.D(_0049_),
    .GATE_N(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[22] ));
 sky130_fd_sc_hd__dlxtn_1 _1978_ (.D(_0050_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[23] ));
 sky130_fd_sc_hd__dlxtn_1 _1979_ (.D(_0051_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[24] ));
 sky130_fd_sc_hd__dlxtn_1 _1980_ (.D(_0052_),
    .GATE_N(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[25] ));
 sky130_fd_sc_hd__dlxtn_1 _1981_ (.D(_0053_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[26] ));
 sky130_fd_sc_hd__dlxtn_1 _1982_ (.D(_0054_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[27] ));
 sky130_fd_sc_hd__dlxtn_1 _1983_ (.D(_0055_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[28] ));
 sky130_fd_sc_hd__dlxtn_1 _1984_ (.D(_0056_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[29] ));
 sky130_fd_sc_hd__dlxtn_1 _1985_ (.D(_0058_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[30] ));
 sky130_fd_sc_hd__dlxtn_1 _1986_ (.D(_0059_),
    .GATE_N(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[31] ));
 sky130_fd_sc_hd__dlxtn_1 _1987_ (.D(_0060_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[32] ));
 sky130_fd_sc_hd__dlxtn_1 _1988_ (.D(_0061_),
    .GATE_N(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tokenflow_inst.i3.ydata[33] ));
 sky130_fd_sc_hd__buf_2 _1989_ (.A(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.ydata[50] ));
 sky130_fd_sc_hd__buf_2 _1990_ (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.ydata[51] ));
 sky130_fd_sc_hd__buf_2 _1991_ (.A(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.ydata[52] ));
 sky130_fd_sc_hd__buf_2 _1992_ (.A(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.ydata[53] ));
 sky130_fd_sc_hd__buf_2 _1993_ (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.ydata[51] ));
 sky130_fd_sc_hd__buf_2 _1994_ (.A(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.ydata[52] ));
 sky130_fd_sc_hd__buf_2 _1995_ (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _1996_ (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _1997_ (.A(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _1998_ (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__buf_2 _1999_ (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__buf_2 _2000_ (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__buf_2 _2001_ (.A(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _2002_ (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__clkbuf_4 _2003_ (.A(\tokenflow_inst.i3.ydata[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _2004_ (.A(\tokenflow_inst.i3.ydata[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__buf_2 _2005_ (.A(\tokenflow_inst.i3.ydata[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _2006_ (.A(\tokenflow_inst.i3.ydata[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__buf_6 _2007_ (.A(\tokenflow_inst.i10.cg.b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i1.c.maj  (.A(_0026_),
    .B(_0027_),
    .C(\tokenflow_inst.i1.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i1.c.q ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i10.cg.maj  (.A(_0028_),
    .B(_0029_),
    .C(\tokenflow_inst.i10.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i10.cg.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i10.d0.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i10.d0.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i10.d0.inv_chain[1] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i11.i.cg.maj  (.A(_0030_),
    .B(_0031_),
    .C(\tokenflow_inst.i11.i.cg.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i11.i.cg.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i11.i.d0.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i11.i.d0.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[1] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i2.cg1.maj  (.A(_0032_),
    .B(_0033_),
    .C(\tokenflow_inst.i2.cg1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i2.cg1.q ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i2.cg2.maj  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .B(_0032_),
    .C(\tokenflow_inst.i2.cg2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i2.cg2.q ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i2.cg3.maj  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .B(_0034_),
    .C(\tokenflow_inst.i2.cg3.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i2.cg3.q ));
 sky130_fd_sc_hd__maj3_4 \tokenflow_inst.i3.cg_elem.maj  (.A(_0115_),
    .B(_0114_),
    .C(\tokenflow_inst.i2.cg2.a ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i2.cg2.a ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i3.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i3.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i3.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[3] ));
 sky130_fd_sc_hd__maj3_2 \tokenflow_inst.i6.cg_elem.maj  (.A(net46),
    .B(_0196_),
    .C(\tokenflow_inst.i6.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[10].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[11] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[11].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[12] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[12].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[13] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[13].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[14] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[14].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[15] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[15].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[16] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[16].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[17] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[17].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[18] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[18].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[19] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[19].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[20] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[20].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[21] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[21].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[22] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[22].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[23] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[23].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[24] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[24].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[25] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[25].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[26] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[26].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[27] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[27].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[28] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[28].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[29] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[29].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[30] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[3] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[30].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[31] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[31].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[32] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[32].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[33] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[33].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[34] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[34].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[35] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[35].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[36] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[36].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[37] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[37].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[38] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[38].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[39] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[39].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[40] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[3].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[4] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[40].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[41] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[41].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[42] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[42].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[43] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[43].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[44] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[44].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[45] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[45].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[46] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[46].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[47] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[47].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[48] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[48].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[49] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[49].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[50] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[4].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[5] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[50].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[51] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[51].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[52] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[5].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[6] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[6].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[7] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[7].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[8] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[8].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[9] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i6.d0_elem.genblk1[9].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[10] ));
 sky130_fd_sc_hd__maj3_4 \tokenflow_inst.i78.cg_elem.maj  (.A(_0273_),
    .B(_0272_),
    .C(\tokenflow_inst.i78.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i78.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i78.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i78.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[3] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i8.cg_elem.maj  (.A(net27),
    .B(_0350_),
    .C(\tokenflow_inst.i8.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[10].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[11] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[11].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[12] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[12].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[13] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[13].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[14] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[14].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[15] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[15].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[16] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[16].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[17] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[17].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[18] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[18].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[19] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[19].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[20] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[20].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[21] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[21].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[22] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[22].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[23] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[23].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[24] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[24].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[25] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[25].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[26] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[26].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[27] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[27].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[28] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[28].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[29] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[29].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[30] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[3] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[30].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[31] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[31].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[32] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[32].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[33] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[33].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[34] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[34].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[35] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[35].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[36] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[36].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[37] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[37].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[38] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[38].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[39] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[39].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[40] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[3].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[4] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[40].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[41] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[41].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[42] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[42].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[43] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[43].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[44] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[44].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[45] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[45].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[46] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[46].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[47] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[47].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[48] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[48].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[49] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[49].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[50] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[4].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[5] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[50].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[51] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[51].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[52] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[5].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[6] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[6].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[7] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[7].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[8] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[8].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[9] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.i8.d0_elem.genblk1[9].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[10] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.i9.c.maj  (.A(_0351_),
    .B(\tokenflow_inst.i10.d0.inv_chain[0] ),
    .C(\tokenflow_inst.i9.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.i9.c.q ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.ii1.cg_elem.maj  (.A(net49),
    .B(_0026_),
    .C(\tokenflow_inst.ii1.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii1.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.ii1.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.ii1.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.ii2.cg_elem.maj  (.A(net56),
    .B(_0381_),
    .C(\tokenflow_inst.ii2.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii2.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.ii2.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.ii2.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.ii2.d0_elem.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[2] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.ii3.i.cg_elem.maj  (.A(_0408_),
    .B(_0409_),
    .C(\tokenflow_inst.ii3.i.cg_elem.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii3.i.cg_elem.q ));
 sky130_fd_sc_hd__clkbuf_1 \tokenflow_inst.ii3.i.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ));
 sky130_fd_sc_hd__maj3_1 \tokenflow_inst.ii4.c.maj  (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .B(_0410_),
    .C(\tokenflow_inst.ii4.c.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tokenflow_inst.ii4.c.q ));
 sky130_fd_sc_hd__conb_1 _1995__137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net137));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_6 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_2 fanout3 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 fanout4 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_2 fanout5 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_2 fanout6 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_2 fanout7 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_2 fanout9 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(_0778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout15 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(_0777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(\tokenflow_inst.i8.ydata[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(\tokenflow_inst.i8.ydata[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout45 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout46 (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_1 fanout49 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_1 fanout56 (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 fanout60 (.A(\tokenflow_inst.i6.ydata[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_1 fanout62 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(\tokenflow_inst.i6.ydata[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_1 fanout72 (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__buf_1 fanout91 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__buf_1 fanout93 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__buf_1 fanout98 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 fanout101 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 fanout104 (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__buf_1 fanout105 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__buf_1 fanout107 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 fanout117 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__buf_1 fanout119 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_1 fanout120 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__buf_8 fanout121 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__buf_1 fanout126 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__buf_8 fanout130 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__conb_1 _1989__131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net131));
 sky130_fd_sc_hd__conb_1 _1990__132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net132));
 sky130_fd_sc_hd__conb_1 _1991__133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net133));
 sky130_fd_sc_hd__conb_1 _1992__134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net134));
 sky130_fd_sc_hd__conb_1 _1993__135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net135));
 sky130_fd_sc_hd__conb_1 _1994__136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net136));
 sky130_fd_sc_hd__conb_1 _1996__138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net138));
 sky130_fd_sc_hd__conb_1 _1997__139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net139));
 sky130_fd_sc_hd__conb_1 _1998__140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net140));
 sky130_fd_sc_hd__conb_1 _1999__141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net141));
 sky130_fd_sc_hd__conb_1 _2000__142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net142));
 sky130_fd_sc_hd__conb_1 _2001__143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net143));
 sky130_fd_sc_hd__conb_1 _2002__144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net144));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_144 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_215 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_131 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_188 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_167 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_83 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_186 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
